
.SUBCKT sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Y C2 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 net62 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net62 C2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_8 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net36 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net36 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net31 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net35 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net31 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Y A net35 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
rI12 VGND LO short
rI11 HI VPWR short
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net118 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net118 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net181 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net181 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net83 net121 net109 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net109 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net102 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net94 M1 net102 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net121 clkneg net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net83 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net82 net83 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net121 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net166 net83 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net83 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net121 clkpos net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net83 net121 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net145 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net145 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net145 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net83 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net121 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net129 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net80 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net129 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net97 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net89 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net89 S1 net97 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net80 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net141 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net141 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net192 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net192 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net156 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net141 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net141 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net128 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net111 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net96 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net88 S1 net96 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net111 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net140 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net140 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net191 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net191 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net168 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net168 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net155 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net140 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net140 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=1 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=5 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=5 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net121 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net121 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net112 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net56 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net112 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net56 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net52 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net52 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net112 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net112 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net107 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net107 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net87 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net87 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net53 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net53 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net44 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net96 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net76 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net76 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net55 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net55 net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 X net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net55 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net55 net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 X net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
MMIN1 Ab X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 net43 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net43 net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 X net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 net43 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net43 net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net56 net48 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net52 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net48 net44 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net44 net52 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net56 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net56 net48 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net48 net44 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net44 net52 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net52 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
MI14 net124 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net124 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net68 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net92 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net92 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net85 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net85 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net68 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Q_N S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net193 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net193 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net148 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net168 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net168 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net161 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net161 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net148 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net141 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net141 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Q_N S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
MI14 net115 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net115 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net59 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net79 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net83 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net83 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net79 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net76 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net76 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net59 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net175 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net175 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net172 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net148 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net148 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net172 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net128 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj31 sndNCINn3 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND A sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR A sndPCINp3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 sndPCINp3 CIN majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj31 sndPCINp3 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
MMIN2 COUT net195 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net123 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb mid2 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Bb mid1 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb mid2 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb mid1 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 CIbb CIb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 CIb CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Ab2 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 Abb2 Ab2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 Ab1 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb2 B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab1 Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb2 Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab1 B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT net195 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM net123 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb mid1 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb mid2 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb mid1 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb mid2 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 CIbb CIb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 CIb CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 Ab2 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 Abb2 Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 Ab1 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb2 Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab1 B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb2 B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab1 Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMIP3 SUM net144 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bbb Bb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CINb1 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CINbb2 CINb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CINb2 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CINbb2 mid2 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CINb2 mid1 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bbb mid2 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CINb1 mid1 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net144 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CINb1 mid2 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CINb1 CIN VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CINbb2 CINb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CINb2 CIN VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CINbb2 mid1 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CINb2 mid2 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bbb mid1 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bbb Bb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
MMIP3 SUM net146 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bb2 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb1 mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb1 mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CIb1 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CIbb2 CIb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CIb2 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb1 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb2 mid2 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb2 mid1 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb2 mid2 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb1 mid1 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net146 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb1 mid2 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb1 mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb1 mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CIb1 CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CIbb2 CIb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CIb2 CI VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb1 B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb2 mid1 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb2 mid2 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bb2 mid1 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bb2 B VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_bleeder_1 SHORT VGND VNB VPB VPWR
MI2 net29 SHORT net25 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net25 SHORT net24 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VPWR SHORT net29 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net24 SHORT net16 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net16 SHORT VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_2 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_4 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_8 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_16 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_1 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_2 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_8 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_16 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_3 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_4 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_6 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_8 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_12 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0n_1 A SLEEP_B VGND VNB VPB VPWR X
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net36 A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 sndA SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 net36 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
MI8 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net36 sleepb VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 sleepb SLEEP VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 sleepb sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 sleepb SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 sndA A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1n_1 A SLEEP_B VGND VNB VPB VPWR X
MI23 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 VPWR net44 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 net56 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA net56 net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 net56 SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net44 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X net44 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net44 net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA A net36 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 VPWR net36 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net36 SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputisolatch_1 D SLEEP_B VGND VNB VPB VPWR Q
MI677 Q s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 sleepneg sleeppos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI674 net39 s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 s0 sleepneg net49 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net49 D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 sleeppos net38 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net38 net39 VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 sleeppos SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 sleeppos SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 sleepneg sleeppos VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
MI662 net86 net39 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 sleepneg net86 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net39 s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 s0 sleeppos net69 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net69 D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_16 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 A SLEEP KAPWR VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA net58 net66 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net58 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab net66 KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net66 SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 net66 net58 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net58 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Ab net66 VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 A VGND VPB VPWRIN VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 A LOWLVPWR VGND VNB VPB VPWR X
MI2 net72 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 cross1 net72 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Ab A LOWLVPWR LOWLVPWR pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 X net60 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 net60 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 cross1 Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net72 A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 X net60 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 net60 cross1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 A LOWLVPWR VGND VPB VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
XI1 net59 LO VGND VNB VPB VPWR / sky130_fd_sc_hd__conb_1
XI6 nor2right invright VGND VNB VPB VPWR / sky130_fd_sc_hd__inv_2
XI7 nor2left invleft VGND VNB VPB VPWR / sky130_fd_sc_hd__inv_2
XI4 nd2right nd2right nor2right VGND VNB VPB VPWR /
+ sky130_fd_sc_hd__nor2_2
XI5 nd2left nd2left nor2left VGND VNB VPB VPWR /
+ sky130_fd_sc_hd__nor2_2
XI2 LO LO nd2right VGND VNB VPB VPWR / sky130_fd_sc_hd__nand2_2
XI3 LO LO nd2left VGND VNB VPB VPWR / sky130_fd_sc_hd__nand2_2
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_2 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_4 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_0 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.7 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__probe_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net29 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net29 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net29 X short
.ENDS




.SUBCKT sky130_fd_sc_hd__probec_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net33 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net33 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net33 X short
rI120 VGND met5vgnd short
rI119 VPWR met5vpwr short
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net153 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net153 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net128 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net128 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net103 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net103 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net87 net153 net117 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net117 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net110 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net98 M1 net110 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net153 clkneg net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net87 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net93 net87 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net153 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net87 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net87 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net153 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net87 net153 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net87 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net153 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net83 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net83 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net159 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net159 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net138 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net199 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net199 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net98 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net98 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI27 net243 S1 net215 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net230 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net227 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net199 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net215 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net206 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net199 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net227 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net230 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net243 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net195 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net195 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net130 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net130 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net107 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI34 S0 clkpos net219 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net239 S1 net187 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net230 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net199 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net230 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net219 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net239 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net199 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net195 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net187 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net195 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net212 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net196 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net212 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net196 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net104 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net104 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net177 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net160 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net177 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net160 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net196 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net189 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net196 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net189 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net138 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net123 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net123 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net235 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net235 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net203 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net203 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net240 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net240 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net180 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net180 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net103 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net103 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net179 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net179 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net135 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net135 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net227 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net227 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net206 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net190 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net190 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net163 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net163 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd2_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_1 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_2 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_4 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_1 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_2 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_4 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS





























































































.subckt user_project_wrapper VGND VPWR wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
XFILLER_100_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09671_ _10761_/A VGND VGND VPWR VPWR _09672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08622_ _08622_/A VGND VGND VPWR VPWR _10112_/B sky130_fd_sc_hd__inv_2
XFILLER_27_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08553_ _09470_/B VGND VGND VPWR VPWR _08688_/A sky130_fd_sc_hd__buf_1
XFILLER_35_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08484_ _08275_/A _08357_/B _08480_/Y _08483_/X VGND VGND VPWR VPWR _08625_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09105_ _08674_/Y _09028_/A _09030_/B VGND VGND VPWR VPWR _09105_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09036_ _09555_/B _09036_/B VGND VGND VPWR VPWR _09037_/B sky130_fd_sc_hd__or2_1
XFILLER_117_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09938_ _09936_/X _09937_/Y _09791_/C _09874_/X _09888_/X VGND VGND VPWR VPWR _09938_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_100_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09869_ _09451_/Y _09868_/X _09472_/X VGND VGND VPWR VPWR _09869_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11900_ _11900_/A VGND VGND VPWR VPWR _11900_/Y sky130_fd_sc_hd__inv_2
X_12880_ _12938_/A VGND VGND VPWR VPWR _14532_/A sky130_fd_sc_hd__buf_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11831_ _12826_/A _11791_/B _11791_/A _11791_/B VGND VGND VPWR VPWR _11831_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14517_/X _14549_/X _14517_/X _14549_/X VGND VGND VPWR VPWR _14582_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13501_/A _13501_/B VGND VGND VPWR VPWR _13501_/Y sky130_fd_sc_hd__nand2_1
X_11762_ _10381_/A _11761_/A _10381_/Y _11805_/B VGND VGND VPWR VPWR _11764_/B sky130_fd_sc_hd__o22a_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _12788_/A VGND VGND VPWR VPWR _13995_/A sky130_fd_sc_hd__buf_1
X_14481_ _14481_/A VGND VGND VPWR VPWR _15196_/A sky130_fd_sc_hd__buf_1
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10713_ _09978_/A _09652_/B _09652_/Y VGND VGND VPWR VPWR _10713_/X sky130_fd_sc_hd__o21a_1
X_16220_ _16253_/B VGND VGND VPWR VPWR _16320_/A sky130_fd_sc_hd__buf_1
X_13432_ _13428_/Y _13430_/Y _13431_/Y VGND VGND VPWR VPWR _13436_/B sky130_fd_sc_hd__o21ai_1
X_10644_ _11907_/A _10644_/B VGND VGND VPWR VPWR _10644_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16151_ _15818_/X _16150_/X _15818_/X _16150_/X VGND VGND VPWR VPWR _16152_/B sky130_fd_sc_hd__a2bb2o_1
X_13363_ _13363_/A _13363_/B VGND VGND VPWR VPWR _13363_/X sky130_fd_sc_hd__or2_1
X_10575_ _13516_/A _10663_/B _13516_/A _10663_/B VGND VGND VPWR VPWR _10575_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12314_ _12322_/A VGND VGND VPWR VPWR _15512_/A sky130_fd_sc_hd__buf_1
X_15102_ _12380_/X _15101_/X _12380_/X _15101_/X VGND VGND VPWR VPWR _15104_/B sky130_fd_sc_hd__a2bb2o_1
Xrebuffer7 rebuffer8/X VGND VGND VPWR VPWR rebuffer7/X sky130_fd_sc_hd__dlygate4sd1_1
X_16082_ _16084_/A _16084_/B VGND VGND VPWR VPWR _16082_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13294_ _14737_/A _13294_/B VGND VGND VPWR VPWR _13294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12245_ _14058_/A _12209_/B _12209_/Y _12244_/X VGND VGND VPWR VPWR _12245_/X sky130_fd_sc_hd__a2bb2o_1
X_15033_ _15076_/A _15031_/X _15032_/X VGND VGND VPWR VPWR _15033_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12176_ _12176_/A VGND VGND VPWR VPWR _12268_/B sky130_fd_sc_hd__inv_2
XFILLER_110_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11127_ _12187_/A VGND VGND VPWR VPWR _13716_/A sky130_fd_sc_hd__buf_1
XFILLER_1_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15935_ _15891_/X _15934_/Y _15891_/X _15934_/Y VGND VGND VPWR VPWR _15954_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11058_ _12232_/A VGND VGND VPWR VPWR _11792_/A sky130_fd_sc_hd__inv_2
XFILLER_37_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15866_ _15866_/A VGND VGND VPWR VPWR _15896_/A sky130_fd_sc_hd__inv_2
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10009_ _10009_/A _10009_/B VGND VGND VPWR VPWR _10035_/B sky130_fd_sc_hd__nor2_1
X_14817_ _14812_/A _14812_/B _14812_/Y _14816_/X VGND VGND VPWR VPWR _14817_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15797_ _15671_/A _15671_/B _15671_/Y VGND VGND VPWR VPWR _15797_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14748_ _14668_/X _14682_/A _14681_/X VGND VGND VPWR VPWR _14748_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14679_ _14670_/X _14678_/X _14670_/X _14678_/X VGND VGND VPWR VPWR _14681_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16418_ _16473_/Q VGND VGND VPWR VPWR _16419_/B sky130_fd_sc_hd__inv_2
XFILLER_32_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16349_ _16335_/X _16348_/Y _16335_/X _16348_/Y VGND VGND VPWR VPWR _16349_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09723_ _09723_/A _09723_/B VGND VGND VPWR VPWR _09723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09654_ _09981_/A _09654_/B VGND VGND VPWR VPWR _09654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08605_ _09250_/A _09217_/B _10015_/A _08604_/Y VGND VGND VPWR VPWR _08605_/X sky130_fd_sc_hd__o22a_1
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09585_ _09993_/A _09662_/B VGND VGND VPWR VPWR _09585_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08536_ _08535_/A _08453_/Y _08535_/Y _08453_/A VGND VGND VPWR VPWR _10119_/B sky130_fd_sc_hd__o22a_1
XFILLER_51_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08467_ _09146_/A VGND VGND VPWR VPWR _08704_/B sky130_fd_sc_hd__inv_2
XFILLER_23_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08398_ _09232_/B VGND VGND VPWR VPWR _08398_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10360_ _13525_/A _10319_/B _10319_/X _10359_/X VGND VGND VPWR VPWR _10360_/X sky130_fd_sc_hd__o22a_1
XFILLER_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10291_ _12706_/A _10291_/B VGND VGND VPWR VPWR _10291_/X sky130_fd_sc_hd__or2_1
X_09019_ _09019_/A VGND VGND VPWR VPWR _09531_/B sky130_fd_sc_hd__inv_2
X_12030_ _13190_/A _12055_/B VGND VGND VPWR VPWR _12030_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13981_ _14836_/A _13981_/B VGND VGND VPWR VPWR _13981_/Y sky130_fd_sc_hd__nor2_1
X_15720_ _14923_/X _15719_/X _14923_/X _15719_/X VGND VGND VPWR VPWR _15721_/B sky130_fd_sc_hd__a2bb2oi_1
X_12932_ _12932_/A _12932_/B VGND VGND VPWR VPWR _12932_/Y sky130_fd_sc_hd__nand2_1
X_15651_ _15651_/A VGND VGND VPWR VPWR _15651_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14602_ _14593_/X _14601_/X _14593_/X _14601_/X VGND VGND VPWR VPWR _14604_/B sky130_fd_sc_hd__a2bb2o_1
X_12863_ _12863_/A _12863_/B VGND VGND VPWR VPWR _12863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15582_ _16051_/A VGND VGND VPWR VPWR _15685_/A sky130_fd_sc_hd__inv_2
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12782_/X _12793_/Y _12782_/X _12793_/Y VGND VGND VPWR VPWR _12858_/B sky130_fd_sc_hd__a2bb2o_1
X_11814_ _12771_/A _11848_/A _11813_/Y VGND VGND VPWR VPWR _11814_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14532_/A _14532_/B _14532_/Y VGND VGND VPWR VPWR _14533_/X sky130_fd_sc_hd__a21o_1
XFILLER_42_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11745_ _11745_/A _11745_/B VGND VGND VPWR VPWR _11745_/X sky130_fd_sc_hd__or2_1
XFILLER_14_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ _14451_/Y _14462_/X _14463_/Y VGND VGND VPWR VPWR _14464_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16203_ _16099_/A _16099_/B _16099_/Y VGND VGND VPWR VPWR _16203_/X sky130_fd_sc_hd__o21a_1
X_13415_ _13357_/X _13414_/X _13357_/X _13414_/X VGND VGND VPWR VPWR _13415_/Y sky130_fd_sc_hd__a2bb2oi_2
X_11676_ _11617_/Y _11621_/Y _12425_/A _11615_/A VGND VGND VPWR VPWR _11676_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_41_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14395_ _15590_/A _14393_/X _14394_/X VGND VGND VPWR VPWR _14395_/X sky130_fd_sc_hd__o21a_1
X_10627_ _13001_/A _10626_/B _10764_/A _10626_/Y VGND VGND VPWR VPWR _10627_/X sky130_fd_sc_hd__o2bb2a_1
X_16134_ _16122_/X _16133_/X _16122_/X _16133_/X VGND VGND VPWR VPWR _16135_/B sky130_fd_sc_hd__a2bb2o_1
X_13346_ _13349_/A VGND VGND VPWR VPWR _15470_/A sky130_fd_sc_hd__buf_1
X_10558_ _10966_/A _11207_/A VGND VGND VPWR VPWR _10559_/A sky130_fd_sc_hd__or2_1
XFILLER_127_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16065_ _16046_/A _16046_/B _16046_/Y VGND VGND VPWR VPWR _16065_/Y sky130_fd_sc_hd__o21ai_1
X_13277_ _13264_/Y _13275_/X _13276_/Y VGND VGND VPWR VPWR _13278_/A sky130_fd_sc_hd__o21ai_1
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12228_ _12228_/A _12137_/X VGND VGND VPWR VPWR _12228_/X sky130_fd_sc_hd__or2b_1
X_10489_ _13625_/A _10531_/B VGND VGND VPWR VPWR _10489_/Y sky130_fd_sc_hd__nor2_1
X_15016_ _15038_/A _15038_/B VGND VGND VPWR VPWR _15067_/A sky130_fd_sc_hd__and2_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12159_ _12158_/Y _12067_/X _12101_/Y VGND VGND VPWR VPWR _12159_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15918_ _15970_/A _15970_/B VGND VGND VPWR VPWR _15918_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15849_ _14184_/A _15848_/X _12633_/X VGND VGND VPWR VPWR _15849_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09370_ _10238_/A VGND VGND VPWR VPWR _09371_/B sky130_fd_sc_hd__buf_1
X_08321_ _08321_/A input19/X VGND VGND VPWR VPWR _08322_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08252_ input17/X VGND VGND VPWR VPWR _08326_/A sky130_fd_sc_hd__inv_2
XFILLER_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09706_ _09689_/A _09689_/B _09692_/A VGND VGND VPWR VPWR _09963_/A sky130_fd_sc_hd__a21bo_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09637_ _09958_/A _09640_/B VGND VGND VPWR VPWR _09637_/Y sky130_fd_sc_hd__nor2_1
X_09568_ _09560_/X _09567_/X _09560_/X _09567_/X VGND VGND VPWR VPWR _09569_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08519_ _09525_/A VGND VGND VPWR VPWR _09476_/B sky130_fd_sc_hd__inv_2
XFILLER_90_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11530_ _11530_/A VGND VGND VPWR VPWR _11530_/Y sky130_fd_sc_hd__inv_2
X_09499_ _08831_/X _09463_/X _08831_/X _09463_/X VGND VGND VPWR VPWR _09500_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11461_ _08983_/X _11460_/X _08983_/X _11460_/X VGND VGND VPWR VPWR _11462_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14180_ _15906_/A _14278_/B VGND VGND VPWR VPWR _14180_/Y sky130_fd_sc_hd__nor2_1
X_11392_ _14103_/A VGND VGND VPWR VPWR _12344_/A sky130_fd_sc_hd__inv_2
X_13200_ _13200_/A _13200_/B VGND VGND VPWR VPWR _13200_/Y sky130_fd_sc_hd__nand2_1
X_10412_ _09297_/Y _10411_/Y _09297_/A _10411_/A _09392_/A VGND VGND VPWR VPWR _12825_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_109_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13131_ _14149_/A VGND VGND VPWR VPWR _13450_/A sky130_fd_sc_hd__buf_1
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10343_ _10352_/A _10342_/X _10352_/A _10342_/X VGND VGND VPWR VPWR _10355_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_124_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13062_ _15246_/A _13117_/B VGND VGND VPWR VPWR _13062_/Y sky130_fd_sc_hd__nor2_1
X_10274_ _11729_/A VGND VGND VPWR VPWR _11724_/A sky130_fd_sc_hd__buf_1
XFILLER_3_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12013_ _11977_/X _12012_/Y _11977_/X _12012_/Y VGND VGND VPWR VPWR _12063_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15703_ _15991_/A _15825_/B VGND VGND VPWR VPWR _15703_/Y sky130_fd_sc_hd__nand2_1
X_13964_ _13989_/A VGND VGND VPWR VPWR _14956_/A sky130_fd_sc_hd__buf_1
XFILLER_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13895_ _14664_/A _13858_/B _13858_/Y VGND VGND VPWR VPWR _13895_/Y sky130_fd_sc_hd__o21ai_1
X_12915_ _12914_/A _12914_/B _12914_/Y VGND VGND VPWR VPWR _12915_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15634_ _15632_/A _15633_/A _15632_/Y _15633_/Y _15571_/A VGND VGND VPWR VPWR _16034_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12846_ _12846_/A _12846_/B VGND VGND VPWR VPWR _12846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _12424_/X _15564_/Y _12424_/X _15564_/Y VGND VGND VPWR VPWR _15565_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _15202_/A _14516_/B VGND VGND VPWR VPWR _14516_/X sky130_fd_sc_hd__or2_1
X_12777_ _12777_/A _12777_/B VGND VGND VPWR VPWR _12777_/Y sky130_fd_sc_hd__nand2_1
X_15496_ _15483_/X _15495_/X _15483_/X _15495_/X VGND VGND VPWR VPWR _15548_/B sky130_fd_sc_hd__a2bb2o_1
X_11728_ _11776_/A _11728_/B VGND VGND VPWR VPWR _11728_/X sky130_fd_sc_hd__or2_1
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11659_ _11657_/X _11659_/B VGND VGND VPWR VPWR _11659_/X sky130_fd_sc_hd__and2b_1
XFILLER_80_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14447_ _14434_/X _14446_/X _14434_/X _14446_/X VGND VGND VPWR VPWR _14465_/B sky130_fd_sc_hd__a2bb2o_1
X_14378_ _14378_/A _14378_/B VGND VGND VPWR VPWR _14378_/Y sky130_fd_sc_hd__nand2_1
X_16117_ _16051_/A _16051_/B _16051_/Y VGND VGND VPWR VPWR _16117_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_115_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13329_ _14733_/A _13288_/B _13288_/Y VGND VGND VPWR VPWR _13329_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16048_ _16051_/A _16051_/B VGND VGND VPWR VPWR _16048_/Y sky130_fd_sc_hd__nor2_1
X_08870_ _08986_/A _08986_/B VGND VGND VPWR VPWR _08870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09422_ _09272_/A _09420_/Y _09421_/Y VGND VGND VPWR VPWR _09424_/B sky130_fd_sc_hd__o21ai_2
XFILLER_80_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09353_ _09353_/A VGND VGND VPWR VPWR _09353_/Y sky130_fd_sc_hd__inv_2
X_08304_ _08304_/A VGND VGND VPWR VPWR _08304_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09284_ _09462_/B _09801_/A _09227_/X VGND VGND VPWR VPWR _09284_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08235_ input7/X _08235_/B VGND VGND VPWR VPWR _08238_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08999_ _11409_/B VGND VGND VPWR VPWR _11391_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10961_ _12080_/A VGND VGND VPWR VPWR _11997_/A sky130_fd_sc_hd__inv_2
X_13680_ _14501_/A _13687_/B VGND VGND VPWR VPWR _13680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12700_ _12700_/A _12700_/B VGND VGND VPWR VPWR _12700_/Y sky130_fd_sc_hd__nor2_1
X_12631_ _12631_/A _12631_/B VGND VGND VPWR VPWR _12631_/X sky130_fd_sc_hd__or2_1
X_10892_ _10892_/A _09407_/X VGND VGND VPWR VPWR _10893_/A sky130_fd_sc_hd__or2b_1
XFILLER_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12562_ _12559_/Y _12561_/Y _12559_/A _12561_/A _12501_/A VGND VGND VPWR VPWR _12625_/B
+ sky130_fd_sc_hd__o221a_1
X_15350_ _15363_/A _15348_/X _15349_/X VGND VGND VPWR VPWR _15350_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14301_ _13444_/A _13444_/B _13444_/Y VGND VGND VPWR VPWR _14301_/X sky130_fd_sc_hd__o21a_1
X_12493_ _12407_/A _12407_/B _12407_/Y _12409_/A VGND VGND VPWR VPWR _12493_/Y sky130_fd_sc_hd__a2bb2oi_1
X_15281_ _14665_/A _15243_/B _15243_/Y _15280_/X VGND VGND VPWR VPWR _15281_/X sky130_fd_sc_hd__a2bb2o_1
X_11513_ _11516_/A VGND VGND VPWR VPWR _11513_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14232_ _12604_/X _14232_/B VGND VGND VPWR VPWR _14232_/X sky130_fd_sc_hd__and2b_1
X_11444_ _11255_/X _11443_/Y _11255_/X _11443_/Y VGND VGND VPWR VPWR _12554_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14163_ _12649_/Y _14163_/B VGND VGND VPWR VPWR _14163_/X sky130_fd_sc_hd__and2b_1
X_11375_ _14058_/A _11197_/B _11197_/Y VGND VGND VPWR VPWR _11375_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14094_ _15464_/A _14036_/B _14036_/A _14036_/B VGND VGND VPWR VPWR _14094_/X sky130_fd_sc_hd__a2bb2o_1
X_13114_ _13072_/Y _13112_/X _13113_/Y VGND VGND VPWR VPWR _13114_/X sky130_fd_sc_hd__o21a_1
X_10326_ _10325_/A _10325_/B _10325_/Y VGND VGND VPWR VPWR _10326_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13045_/A _13032_/X VGND VGND VPWR VPWR _13045_/X sky130_fd_sc_hd__or2b_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _09275_/B _10244_/B _10244_/X _10569_/A VGND VGND VPWR VPWR _10688_/A sky130_fd_sc_hd__a22o_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10188_ _10242_/B _10155_/B _10155_/Y _10819_/A VGND VGND VPWR VPWR _10973_/A sky130_fd_sc_hd__o2bb2a_1
X_14996_ _14996_/A _15728_/A VGND VGND VPWR VPWR _16125_/A sky130_fd_sc_hd__or2_1
XFILLER_66_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13947_ _13921_/Y _13945_/X _13946_/Y VGND VGND VPWR VPWR _13947_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15617_ _15617_/A VGND VGND VPWR VPWR _15617_/Y sky130_fd_sc_hd__inv_2
X_13878_ _13866_/X _13877_/Y _13866_/X _13877_/Y VGND VGND VPWR VPWR _13981_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12829_ _12829_/A _12829_/B VGND VGND VPWR VPWR _12829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15548_ _15548_/A _15548_/B VGND VGND VPWR VPWR _15579_/B sky130_fd_sc_hd__or2_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15479_ _14798_/A _15458_/B _15458_/Y _15478_/X VGND VGND VPWR VPWR _15479_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_30_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09971_ _09971_/A VGND VGND VPWR VPWR _09971_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08922_ _08922_/A _08922_/B VGND VGND VPWR VPWR _09293_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08853_ _08916_/A _08913_/B VGND VGND VPWR VPWR _08937_/B sky130_fd_sc_hd__or2_1
XFILLER_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08784_ _08786_/B VGND VGND VPWR VPWR _08784_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09405_ _09403_/X _09101_/A _08664_/X _09404_/Y VGND VGND VPWR VPWR _09407_/B sky130_fd_sc_hd__o22a_1
XFILLER_111_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09336_ _08778_/A _08776_/Y _10041_/A _09335_/X VGND VGND VPWR VPWR _09336_/X sky130_fd_sc_hd__o22a_1
X_09267_ _09259_/X _08899_/Y _09259_/X _08899_/Y VGND VGND VPWR VPWR _10243_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09198_ _09198_/A VGND VGND VPWR VPWR _09198_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11160_ _13504_/A _11304_/B _13504_/A _11304_/B VGND VGND VPWR VPWR _11160_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11091_ _13902_/A _11091_/B VGND VGND VPWR VPWR _11091_/X sky130_fd_sc_hd__or2_1
X_10111_ _10111_/A _10111_/B VGND VGND VPWR VPWR _10112_/A sky130_fd_sc_hd__or2_1
XFILLER_88_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10042_ _10027_/X _10041_/Y _10027_/X _10041_/Y VGND VGND VPWR VPWR _10083_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14850_ _14835_/X _14849_/X _14835_/X _14849_/X VGND VGND VPWR VPWR _14953_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14781_ _14738_/X _14780_/X _14738_/X _14780_/X VGND VGND VPWR VPWR _14782_/B sky130_fd_sc_hd__a2bb2o_1
X_13801_ _13801_/A _13775_/X VGND VGND VPWR VPWR _13801_/X sky130_fd_sc_hd__or2b_1
XFILLER_63_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13732_ _13769_/A _13769_/B VGND VGND VPWR VPWR _13810_/A sky130_fd_sc_hd__and2_1
X_11993_ _10678_/A _11922_/A _10811_/B _11992_/Y VGND VGND VPWR VPWR _11994_/A sky130_fd_sc_hd__o22a_1
XFILLER_29_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10944_ _13641_/A _10944_/B VGND VGND VPWR VPWR _10944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16451_ _16437_/D _16419_/B _16445_/X _16448_/X VGND VGND VPWR VPWR _16451_/X sky130_fd_sc_hd__o211a_1
X_10875_ _10875_/A _10875_/B VGND VGND VPWR VPWR _10875_/X sky130_fd_sc_hd__and2_1
X_13663_ _13632_/A _13662_/Y _13632_/A _13662_/Y VGND VGND VPWR VPWR _13697_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16382_ _16312_/Y _16381_/Y _16312_/Y _16381_/Y VGND VGND VPWR VPWR _16396_/C sky130_fd_sc_hd__a2bb2o_1
X_12614_ _12610_/Y _12613_/Y _12610_/A _12613_/A _12499_/A VGND VGND VPWR VPWR _14235_/B
+ sky130_fd_sc_hd__o221a_1
X_15402_ _15402_/A _15402_/B VGND VGND VPWR VPWR _15402_/X sky130_fd_sc_hd__or2_1
X_13594_ _13556_/A _13556_/B _13557_/A VGND VGND VPWR VPWR _13594_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12545_ _15540_/A VGND VGND VPWR VPWR _14916_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15333_ _15333_/A _15333_/B VGND VGND VPWR VPWR _15333_/X sky130_fd_sc_hd__or2_1
XFILLER_61_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12476_ _13463_/A _12478_/B VGND VGND VPWR VPWR _12476_/Y sky130_fd_sc_hd__nor2_1
X_15264_ _15264_/A _15264_/B VGND VGND VPWR VPWR _15264_/Y sky130_fd_sc_hd__nand2_1
X_14215_ _12622_/X _14214_/X _12622_/X _14214_/X VGND VGND VPWR VPWR _14260_/B sky130_fd_sc_hd__a2bb2o_1
X_11427_ _13341_/A _11236_/B _11236_/Y VGND VGND VPWR VPWR _11427_/Y sky130_fd_sc_hd__o21ai_1
X_15195_ _15152_/X _15194_/Y _15152_/X _15194_/Y VGND VGND VPWR VPWR _15196_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14146_ _14140_/X _14143_/Y _14408_/A _14145_/Y VGND VGND VPWR VPWR _14146_/X sky130_fd_sc_hd__o22a_1
XFILLER_4_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11358_ _08979_/X _11357_/X _08979_/X _11357_/X VGND VGND VPWR VPWR _11359_/B sky130_fd_sc_hd__a2bb2oi_2
X_10309_ _10309_/A _10309_/B VGND VGND VPWR VPWR _10309_/Y sky130_fd_sc_hd__nor2_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14077_ _14077_/A _14056_/X VGND VGND VPWR VPWR _14077_/X sky130_fd_sc_hd__or2b_1
X_11289_ _11289_/A VGND VGND VPWR VPWR _11289_/Y sky130_fd_sc_hd__inv_2
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _14592_/A _13028_/B VGND VGND VPWR VPWR _13028_/X sky130_fd_sc_hd__or2_1
XFILLER_67_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer17 rebuffer18/X VGND VGND VPWR VPWR rebuffer17/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer28 _16318_/A VGND VGND VPWR VPWR _16378_/A1 sky130_fd_sc_hd__dlygate4sd1_1
X_14979_ _14977_/Y _14978_/X _14977_/Y _14978_/X VGND VGND VPWR VPWR _14979_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09121_ _09549_/B _09033_/B _09034_/B VGND VGND VPWR VPWR _09122_/A sky130_fd_sc_hd__a21bo_1
XFILLER_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09052_ _09052_/A VGND VGND VPWR VPWR _09052_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09954_ _09954_/A VGND VGND VPWR VPWR _09954_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _09885_/A _09885_/B VGND VGND VPWR VPWR _09886_/B sky130_fd_sc_hd__or2_1
X_08905_ _08904_/X _08810_/B _08810_/Y VGND VGND VPWR VPWR _08905_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _10018_/A _10124_/A VGND VGND VPWR VPWR _08836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08767_ _10132_/A VGND VGND VPWR VPWR _08770_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08698_ _10008_/A VGND VGND VPWR VPWR _09478_/A sky130_fd_sc_hd__buf_1
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10660_ _10660_/A _10660_/B VGND VGND VPWR VPWR _10660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09319_ _08572_/A _09858_/A _09318_/Y _09244_/X VGND VGND VPWR VPWR _09319_/X sky130_fd_sc_hd__o22a_1
X_10591_ _09971_/Y _10590_/A _09971_/A _10590_/Y _09797_/A VGND VGND VPWR VPWR _11901_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12330_ _12590_/A _12589_/A _12329_/X VGND VGND VPWR VPWR _12334_/B sky130_fd_sc_hd__o21ai_1
XFILLER_107_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12261_ _12261_/A _12261_/B VGND VGND VPWR VPWR _12261_/X sky130_fd_sc_hd__or2_1
XFILLER_5_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11212_ _11449_/A _11212_/B VGND VGND VPWR VPWR _11212_/Y sky130_fd_sc_hd__nand2_1
X_14000_ _13986_/A _13987_/X _13985_/X VGND VGND VPWR VPWR _14000_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12192_ _12255_/A _12191_/Y _12255_/A _12191_/Y VGND VGND VPWR VPWR _12252_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11143_ _10082_/X _11142_/X _10082_/X _11142_/X VGND VGND VPWR VPWR _11144_/B sky130_fd_sc_hd__a2bb2o_1
X_15951_ _16020_/A _15949_/X _15950_/X VGND VGND VPWR VPWR _15951_/X sky130_fd_sc_hd__o21a_1
X_11074_ _13936_/A _12232_/B _11072_/X _11246_/A VGND VGND VPWR VPWR _11074_/X sky130_fd_sc_hd__a31o_1
XFILLER_95_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15882_ _14232_/X _15840_/A _14232_/X _15840_/A VGND VGND VPWR VPWR _15886_/B sky130_fd_sc_hd__a2bb2o_1
X_14902_ _14815_/A _14815_/B _14815_/Y VGND VGND VPWR VPWR _14902_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10025_ _09492_/A _09249_/B _10050_/B _10024_/X VGND VGND VPWR VPWR _10025_/X sky130_fd_sc_hd__o22a_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14833_ _14833_/A _14833_/B VGND VGND VPWR VPWR _14833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14764_ _14833_/A _14833_/B VGND VGND VPWR VPWR _14764_/Y sky130_fd_sc_hd__nand2_1
X_11976_ _13063_/A _11976_/B VGND VGND VPWR VPWR _11976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14695_ _14659_/X _14694_/Y _14659_/X _14694_/Y VGND VGND VPWR VPWR _14737_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13715_ _13710_/X _13714_/Y _13710_/X _13714_/Y VGND VGND VPWR VPWR _13779_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10927_ _09323_/A _10925_/A _09328_/A _10925_/Y _11583_/A VGND VGND VPWR VPWR _12104_/A
+ sky130_fd_sc_hd__a221o_2
X_16434_ _16434_/A _16434_/B VGND VGND VPWR VPWR _16434_/Y sky130_fd_sc_hd__nor2_1
X_13646_ _12852_/A _13584_/B _13645_/Y _13581_/X VGND VGND VPWR VPWR _13646_/X sky130_fd_sc_hd__o22a_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10858_ _10774_/X _10857_/Y _10774_/X _10857_/Y VGND VGND VPWR VPWR _10916_/B sky130_fd_sc_hd__o2bb2a_1
X_16365_ _16357_/X _16464_/Q _16358_/X _16407_/C _16361_/X VGND VGND VPWR VPWR _16464_/D
+ sky130_fd_sc_hd__o221a_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10789_ _13637_/A _10789_/B VGND VGND VPWR VPWR _10789_/Y sky130_fd_sc_hd__nor2_1
X_13577_ _12842_/A _13564_/B _13565_/Y _13576_/X VGND VGND VPWR VPWR _13577_/X sky130_fd_sc_hd__o22a_1
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16296_ _16328_/A _16328_/B VGND VGND VPWR VPWR _16296_/Y sky130_fd_sc_hd__nor2_1
X_12528_ _14120_/A VGND VGND VPWR VPWR _13440_/A sky130_fd_sc_hd__buf_1
X_15316_ _15275_/X _15315_/Y _15275_/X _15315_/Y VGND VGND VPWR VPWR _15337_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12459_ _12458_/Y _12361_/Y _12393_/Y VGND VGND VPWR VPWR _12459_/X sky130_fd_sc_hd__o21a_1
X_15247_ _15193_/A _15193_/B _15193_/Y VGND VGND VPWR VPWR _15247_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15178_ _15178_/A _15178_/B VGND VGND VPWR VPWR _15178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14129_ _14129_/A _14062_/X VGND VGND VPWR VPWR _14129_/X sky130_fd_sc_hd__or2b_1
XFILLER_113_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09670_ _09523_/X _09669_/X _09523_/X _09669_/X VGND VGND VPWR VPWR _10761_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_67_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08621_ _08717_/B VGND VGND VPWR VPWR _08623_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08552_ _09531_/A VGND VGND VPWR VPWR _09470_/B sky130_fd_sc_hd__inv_2
XFILLER_35_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08483_ _08276_/Y _08279_/B _08482_/X VGND VGND VPWR VPWR _08483_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09104_ _09407_/A _09104_/B VGND VGND VPWR VPWR _09104_/X sky130_fd_sc_hd__and2_1
X_09035_ _09553_/B _09035_/B VGND VGND VPWR VPWR _09036_/B sky130_fd_sc_hd__or2_1
XFILLER_117_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09937_ _09937_/A _09937_/B VGND VGND VPWR VPWR _09937_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09868_ _09452_/Y _09867_/X _09470_/X VGND VGND VPWR VPWR _09868_/X sky130_fd_sc_hd__o21a_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09799_ _09799_/A _09799_/B VGND VGND VPWR VPWR _09834_/A sky130_fd_sc_hd__or2_1
X_08819_ _08819_/A _10126_/A VGND VGND VPWR VPWR _08819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11830_ _15143_/A _11835_/B VGND VGND VPWR VPWR _11830_/Y sky130_fd_sc_hd__nor2_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11761_/A VGND VGND VPWR VPWR _11805_/B sky130_fd_sc_hd__inv_2
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10712_ _11942_/A _10712_/B VGND VGND VPWR VPWR _10712_/Y sky130_fd_sc_hd__nand2_1
X_13500_ _11332_/X _13491_/X _11332_/X _13491_/X VGND VGND VPWR VPWR _13501_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _15193_/A _14522_/B VGND VGND VPWR VPWR _14541_/A sky130_fd_sc_hd__and2_1
XFILLER_41_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11692_ _11609_/Y _11689_/Y _11691_/X VGND VGND VPWR VPWR _11692_/Y sky130_fd_sc_hd__o21ai_2
X_13431_ _14106_/A _13431_/B VGND VGND VPWR VPWR _13431_/Y sky130_fd_sc_hd__nand2_1
X_10643_ _10643_/A VGND VGND VPWR VPWR _10643_/Y sky130_fd_sc_hd__inv_2
X_16150_ _15718_/X _16150_/B VGND VGND VPWR VPWR _16150_/X sky130_fd_sc_hd__and2b_1
X_13362_ _13331_/A _13331_/B _13331_/X _13361_/X VGND VGND VPWR VPWR _13362_/X sky130_fd_sc_hd__o22a_1
X_10574_ _10553_/X _10573_/X _10553_/X _10573_/X VGND VGND VPWR VPWR _10663_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16081_ _16028_/X _16080_/X _16028_/X _16080_/X VGND VGND VPWR VPWR _16084_/B sky130_fd_sc_hd__a2bb2o_1
X_12313_ _14084_/A VGND VGND VPWR VPWR _12322_/A sky130_fd_sc_hd__inv_2
X_15101_ _12274_/A _15048_/X _12273_/X VGND VGND VPWR VPWR _15101_/X sky130_fd_sc_hd__o21a_1
Xrebuffer8 rebuffer9/X VGND VGND VPWR VPWR rebuffer8/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13293_ _13293_/A VGND VGND VPWR VPWR _13293_/Y sky130_fd_sc_hd__inv_2
X_15032_ _15032_/A _15032_/B VGND VGND VPWR VPWR _15032_/X sky130_fd_sc_hd__or2_1
XFILLER_123_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12244_ _14056_/A _12212_/B _12212_/Y _12243_/X VGND VGND VPWR VPWR _12244_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12175_ _10970_/A _12084_/A _11140_/B _12174_/Y VGND VGND VPWR VPWR _12176_/A sky130_fd_sc_hd__o22a_1
X_11126_ _12942_/A VGND VGND VPWR VPWR _12187_/A sky130_fd_sc_hd__inv_2
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15934_ _15892_/A _15892_/B _15892_/Y VGND VGND VPWR VPWR _15934_/Y sky130_fd_sc_hd__o21ai_1
X_11057_ _12137_/A _11076_/B VGND VGND VPWR VPWR _11240_/A sky130_fd_sc_hd__and2_1
XFILLER_49_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15865_ _15898_/A _15898_/B VGND VGND VPWR VPWR _15865_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10008_ _10008_/A _10008_/B VGND VGND VPWR VPWR _10008_/X sky130_fd_sc_hd__or2_1
X_14816_ _14815_/A _14815_/B _14047_/X _14815_/Y VGND VGND VPWR VPWR _14816_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_91_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15796_ _15799_/A _15800_/B VGND VGND VPWR VPWR _15796_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14747_ _14666_/X _14746_/Y _14684_/Y VGND VGND VPWR VPWR _14747_/X sky130_fd_sc_hd__o21a_1
X_11959_ _11959_/A VGND VGND VPWR VPWR _11959_/X sky130_fd_sc_hd__buf_1
XFILLER_60_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14678_ _14677_/A _14677_/B _14677_/Y VGND VGND VPWR VPWR _14678_/X sky130_fd_sc_hd__a21o_1
X_16417_ _16466_/Q VGND VGND VPWR VPWR _16437_/B sky130_fd_sc_hd__inv_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13629_ _13629_/A VGND VGND VPWR VPWR _15131_/A sky130_fd_sc_hd__buf_1
XFILLER_20_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16348_ _16336_/A _16336_/B _16336_/Y VGND VGND VPWR VPWR _16348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16279_ _16273_/A _16338_/A _16273_/Y VGND VGND VPWR VPWR _16279_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09722_ _09723_/A _09723_/B VGND VGND VPWR VPWR _09722_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09653_ _09615_/Y _09651_/X _09652_/Y VGND VGND VPWR VPWR _09653_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08604_ _09217_/B VGND VGND VPWR VPWR _08604_/Y sky130_fd_sc_hd__inv_2
X_09584_ _09557_/X _09583_/X _09557_/X _09583_/X VGND VGND VPWR VPWR _09662_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _08535_/A VGND VGND VPWR VPWR _08535_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08466_ _08465_/A _08239_/Y _08465_/Y _08239_/A _08441_/X VGND VGND VPWR VPWR _09146_/A
+ sky130_fd_sc_hd__o221a_2
X_08397_ _08399_/B _08392_/A _08282_/A _08392_/Y _08663_/B VGND VGND VPWR VPWR _09232_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10290_ _13479_/A _10286_/B _10289_/X VGND VGND VPWR VPWR _10291_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09018_ _08778_/A _09014_/Y _09014_/Y _08558_/Y VGND VGND VPWR VPWR _09019_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13980_ _13980_/A _13979_/X VGND VGND VPWR VPWR _13980_/X sky130_fd_sc_hd__or2b_1
XFILLER_58_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12931_ _12899_/Y _12929_/X _12930_/Y VGND VGND VPWR VPWR _12931_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15650_ _15650_/A VGND VGND VPWR VPWR _15650_/Y sky130_fd_sc_hd__inv_2
X_12862_ _12789_/X _12861_/X _12789_/X _12861_/X VGND VGND VPWR VPWR _12863_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14601_ _14600_/A _14600_/B _14600_/Y VGND VGND VPWR VPWR _14601_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11813_ _12771_/A _11848_/A VGND VGND VPWR VPWR _11813_/Y sky130_fd_sc_hd__nor2_1
X_15581_ _15700_/A _15581_/B VGND VGND VPWR VPWR _16051_/A sky130_fd_sc_hd__or2_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12793_ _12783_/A _12783_/B _12783_/Y VGND VGND VPWR VPWR _12793_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14532_/A _14532_/B VGND VGND VPWR VPWR _14532_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11744_ _11742_/A _11742_/B _11742_/X _11743_/Y VGND VGND VPWR VPWR _11757_/B sky130_fd_sc_hd__a22o_1
XFILLER_14_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14463_/A _14463_/B VGND VGND VPWR VPWR _14463_/Y sky130_fd_sc_hd__nand2_1
X_11675_ _12679_/A VGND VGND VPWR VPWR _12425_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16202_ _16257_/A _16258_/B VGND VGND VPWR VPWR _16202_/Y sky130_fd_sc_hd__nor2_1
X_13414_ _15467_/A _13345_/B _13345_/Y VGND VGND VPWR VPWR _13414_/X sky130_fd_sc_hd__a21o_1
X_10626_ _11889_/A _10626_/B VGND VGND VPWR VPWR _10626_/Y sky130_fd_sc_hd__nor2_1
X_16133_ _16061_/X _16133_/B VGND VGND VPWR VPWR _16133_/X sky130_fd_sc_hd__and2b_1
X_14394_ _15964_/A _14394_/B VGND VGND VPWR VPWR _14394_/X sky130_fd_sc_hd__or2_1
X_13345_ _14039_/A _13345_/B VGND VGND VPWR VPWR _13345_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10557_ _09088_/A _10556_/X _09088_/A _10556_/X VGND VGND VPWR VPWR _11207_/A sky130_fd_sc_hd__a2bb2o_2
X_16064_ _16121_/A _16121_/B VGND VGND VPWR VPWR _16138_/A sky130_fd_sc_hd__and2_1
XFILLER_115_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13276_ _14725_/A _13276_/B VGND VGND VPWR VPWR _13276_/Y sky130_fd_sc_hd__nand2_1
X_10488_ _10435_/X _10487_/X _10435_/X _10487_/X VGND VGND VPWR VPWR _10531_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12227_ _12227_/A _12227_/B VGND VGND VPWR VPWR _12227_/Y sky130_fd_sc_hd__nand2_1
X_15015_ _11860_/X _15002_/X _11860_/X _15002_/X VGND VGND VPWR VPWR _15038_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12158_ _12158_/A _12158_/B VGND VGND VPWR VPWR _12158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11109_ _11276_/A VGND VGND VPWR VPWR _14664_/A sky130_fd_sc_hd__buf_1
XFILLER_68_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12089_ _12172_/B _12088_/X _12172_/B _12088_/X VGND VGND VPWR VPWR _12168_/A sky130_fd_sc_hd__a2bb2o_1
X_15917_ _15907_/X _15916_/Y _15907_/X _15916_/Y VGND VGND VPWR VPWR _15970_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15848_ _14190_/A _15847_/X _12631_/X VGND VGND VPWR VPWR _15848_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15779_ _14364_/A _15774_/A _14376_/A VGND VGND VPWR VPWR _16028_/B sky130_fd_sc_hd__a21bo_1
XFILLER_52_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08320_ _08318_/Y _08319_/A _08318_/A _08319_/Y _08304_/X VGND VGND VPWR VPWR _08543_/B
+ sky130_fd_sc_hd__o221a_1
X_08251_ input3/X _08251_/B VGND VGND VPWR VPWR _08322_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09705_ _09705_/A VGND VGND VPWR VPWR _09720_/A sky130_fd_sc_hd__inv_2
XFILLER_74_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09636_ _09952_/A _09631_/B _09632_/Y _09635_/Y VGND VGND VPWR VPWR _09640_/B sky130_fd_sc_hd__o22a_1
XFILLER_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09567_ _09567_/A _09567_/B VGND VGND VPWR VPWR _09567_/X sky130_fd_sc_hd__or2_1
X_08518_ _08701_/A _08518_/B VGND VGND VPWR VPWR _09525_/A sky130_fd_sc_hd__or2_2
X_09498_ _09498_/A _09498_/B VGND VGND VPWR VPWR _09498_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08449_ _08543_/A VGND VGND VPWR VPWR _10010_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11460_ _08875_/X _11460_/B VGND VGND VPWR VPWR _11460_/X sky130_fd_sc_hd__and2b_1
X_11391_ _11391_/A _11391_/B VGND VGND VPWR VPWR _14103_/A sky130_fd_sc_hd__or2_1
X_10411_ _10411_/A VGND VGND VPWR VPWR _10411_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13130_ _13128_/Y _13129_/X _13128_/Y _13129_/X VGND VGND VPWR VPWR _13130_/X sky130_fd_sc_hd__o2bb2a_1
X_10342_ _13479_/A _10286_/B _10289_/A VGND VGND VPWR VPWR _10342_/X sky130_fd_sc_hd__o21ba_1
XFILLER_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13061_ _13025_/X _13060_/X _13025_/X _13060_/X VGND VGND VPWR VPWR _13117_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12012_ _13058_/A _12066_/B _12011_/Y VGND VGND VPWR VPWR _12012_/Y sky130_fd_sc_hd__o21ai_1
X_10273_ _10108_/Y _10272_/Y _10108_/A _10272_/A _10472_/A VGND VGND VPWR VPWR _11729_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15702_ _14404_/X _15701_/Y _14404_/X _15701_/Y VGND VGND VPWR VPWR _15825_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13963_ _13889_/Y _13961_/X _13962_/Y VGND VGND VPWR VPWR _13963_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13894_ _13894_/A VGND VGND VPWR VPWR _15416_/A sky130_fd_sc_hd__buf_1
X_12914_ _12914_/A _12914_/B VGND VGND VPWR VPWR _12914_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15633_ _15633_/A VGND VGND VPWR VPWR _15633_/Y sky130_fd_sc_hd__inv_2
X_12845_ _12816_/Y _12843_/X _12844_/Y VGND VGND VPWR VPWR _12845_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15564_ _15563_/Y _15486_/X _15433_/Y VGND VGND VPWR VPWR _15564_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12776_ _12741_/Y _12774_/X _12775_/Y VGND VGND VPWR VPWR _12776_/X sky130_fd_sc_hd__o21a_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _14557_/A _14513_/X _14514_/X VGND VGND VPWR VPWR _14515_/X sky130_fd_sc_hd__o21a_1
X_11727_ _11783_/A _11719_/B _11719_/Y _11784_/B VGND VGND VPWR VPWR _11728_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15495_ _15443_/A _15443_/B _15443_/A _15443_/B VGND VGND VPWR VPWR _15495_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11658_ _12788_/A _11658_/B VGND VGND VPWR VPWR _11659_/B sky130_fd_sc_hd__or2_1
X_14446_ _14423_/A _14423_/B _14423_/Y VGND VGND VPWR VPWR _14446_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14377_ _15662_/B _14375_/Y _15661_/A VGND VGND VPWR VPWR _14377_/X sky130_fd_sc_hd__o21a_1
X_11589_ _09789_/X _11588_/Y _09789_/X _11588_/Y VGND VGND VPWR VPWR _11590_/B sky130_fd_sc_hd__a2bb2oi_1
X_10609_ _09954_/Y _10608_/A _09954_/A _10608_/Y _09797_/A VGND VGND VPWR VPWR _10628_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16116_ _16119_/A _16119_/B VGND VGND VPWR VPWR _16116_/Y sky130_fd_sc_hd__nor2_1
X_13328_ _13363_/A _13363_/B VGND VGND VPWR VPWR _13391_/A sky130_fd_sc_hd__and2_1
XFILLER_6_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16047_ _16001_/Y _16045_/X _16046_/Y VGND VGND VPWR VPWR _16051_/B sky130_fd_sc_hd__o21ai_2
XFILLER_115_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13259_ _13187_/X _13258_/Y _13187_/X _13258_/Y VGND VGND VPWR VPWR _13279_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09421_ _09421_/A _09421_/B VGND VGND VPWR VPWR _09421_/Y sky130_fd_sc_hd__nand2_1
X_09352_ _09529_/A _09740_/A VGND VGND VPWR VPWR _09353_/A sky130_fd_sc_hd__or2_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08303_ _08303_/A VGND VGND VPWR VPWR _08304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09283_ _10250_/A VGND VGND VPWR VPWR _10252_/A sky130_fd_sc_hd__buf_1
X_08234_ input23/X VGND VGND VPWR VPWR _08235_/B sky130_fd_sc_hd__inv_2
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08998_ _12605_/B VGND VGND VPWR VPWR _11409_/B sky130_fd_sc_hd__inv_2
XFILLER_87_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10960_ _10962_/A VGND VGND VPWR VPWR _10960_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10891_ _12037_/A _10891_/B VGND VGND VPWR VPWR _10891_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09619_ _09500_/A _09500_/B _09500_/Y VGND VGND VPWR VPWR _09619_/X sky130_fd_sc_hd__a21o_1
X_12630_ _14196_/A _12628_/X _12629_/X VGND VGND VPWR VPWR _12630_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12561_ _12561_/A VGND VGND VPWR VPWR _12561_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14300_ _14309_/A _14300_/B VGND VGND VPWR VPWR _15970_/A sky130_fd_sc_hd__nor2_1
X_12492_ _12494_/A _12494_/B VGND VGND VPWR VPWR _12492_/Y sky130_fd_sc_hd__nor2_1
X_15280_ _14588_/A _15246_/B _15246_/Y _15279_/X VGND VGND VPWR VPWR _15280_/X sky130_fd_sc_hd__a2bb2o_1
X_11512_ _11626_/A VGND VGND VPWR VPWR _13496_/A sky130_fd_sc_hd__buf_1
XFILLER_12_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14231_ _14231_/A _14231_/B VGND VGND VPWR VPWR _15881_/A sky130_fd_sc_hd__or2_1
X_11443_ _14028_/A _11218_/B _11218_/Y VGND VGND VPWR VPWR _11443_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14162_ _14282_/A _14162_/B VGND VGND VPWR VPWR _15974_/A sky130_fd_sc_hd__or2_1
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11374_ _12309_/A VGND VGND VPWR VPWR _14120_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13113_ _15252_/A _13113_/B VGND VGND VPWR VPWR _13113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14093_ _14093_/A _14096_/B VGND VGND VPWR VPWR _14093_/Y sky130_fd_sc_hd__nor2_1
X_10325_ _10325_/A _10325_/B VGND VGND VPWR VPWR _10325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13044_ _15237_/A VGND VGND VPWR VPWR _14833_/A sky130_fd_sc_hd__buf_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ _09313_/A _10254_/B _10255_/Y _10469_/A VGND VGND VPWR VPWR _10569_/A sky130_fd_sc_hd__o22a_1
XFILLER_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10187_ _10243_/B _10159_/B _10159_/Y _10681_/A VGND VGND VPWR VPWR _10819_/A sky130_fd_sc_hd__o2bb2a_1
X_14995_ _15752_/A VGND VGND VPWR VPWR _15728_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13946_ _15404_/A _13946_/B VGND VGND VPWR VPWR _13946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15616_ _15616_/A VGND VGND VPWR VPWR _15616_/Y sky130_fd_sc_hd__inv_2
X_13877_ _15110_/A _13975_/B _13876_/Y VGND VGND VPWR VPWR _13877_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12828_ _10620_/A _11716_/A _10521_/A _11717_/B VGND VGND VPWR VPWR _12829_/B sky130_fd_sc_hd__o22a_1
X_15547_ _15500_/X _15545_/X _15586_/B VGND VGND VPWR VPWR _15547_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12759_ _12708_/X _12758_/X _12708_/X _12758_/X VGND VGND VPWR VPWR _12763_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15478_ _14802_/A _15461_/B _15461_/Y _15477_/X VGND VGND VPWR VPWR _15478_/X sky130_fd_sc_hd__a2bb2o_1
X_14429_ _14429_/A _14429_/B VGND VGND VPWR VPWR _14429_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09970_ _09970_/A VGND VGND VPWR VPWR _09970_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08921_ _08930_/A _09101_/A VGND VGND VPWR VPWR _08922_/B sky130_fd_sc_hd__or2_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08852_ _08852_/A _08856_/B VGND VGND VPWR VPWR _08913_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08783_ _10130_/A VGND VGND VPWR VPWR _08786_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09404_ _09404_/A VGND VGND VPWR VPWR _09404_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09335_ _09470_/A _08784_/Y _10044_/A _09325_/X VGND VGND VPWR VPWR _09335_/X sky130_fd_sc_hd__o22a_1
X_09266_ _09266_/A VGND VGND VPWR VPWR _09269_/A sky130_fd_sc_hd__inv_2
XFILLER_21_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09197_ _09146_/X _09150_/S _08505_/B VGND VGND VPWR VPWR _09199_/A sky130_fd_sc_hd__o21ba_1
XFILLER_119_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11090_ _11204_/A _11088_/X _11089_/X VGND VGND VPWR VPWR _11090_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10110_ _10110_/A _10110_/B VGND VGND VPWR VPWR _10111_/A sky130_fd_sc_hd__or2_1
X_10041_ _10041_/A _10041_/B VGND VGND VPWR VPWR _10041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14780_ _14780_/A _14739_/X VGND VGND VPWR VPWR _14780_/X sky130_fd_sc_hd__or2b_1
X_13800_ _14745_/A _13860_/B VGND VGND VPWR VPWR _13800_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11992_ _11992_/A _11992_/B VGND VGND VPWR VPWR _11992_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13731_ _13698_/X _13730_/X _13698_/X _13730_/X VGND VGND VPWR VPWR _13769_/B sky130_fd_sc_hd__a2bb2o_1
X_10943_ _12005_/A VGND VGND VPWR VPWR _13641_/A sky130_fd_sc_hd__buf_1
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16450_ _16445_/X _16448_/X _16474_/Q _16449_/X VGND VGND VPWR VPWR _16450_/X sky130_fd_sc_hd__o22a_1
X_10874_ _10772_/X _10873_/Y _10772_/X _10873_/Y VGND VGND VPWR VPWR _10875_/B sky130_fd_sc_hd__o2bb2a_1
X_13662_ _15128_/A _13634_/B _13634_/Y VGND VGND VPWR VPWR _13662_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16381_ _16381_/A1 _16316_/B _16316_/Y VGND VGND VPWR VPWR _16381_/Y sky130_fd_sc_hd__o21ai_1
X_12613_ _12613_/A VGND VGND VPWR VPWR _12613_/Y sky130_fd_sc_hd__inv_2
X_15401_ _15465_/A _15399_/X _15400_/X VGND VGND VPWR VPWR _15401_/X sky130_fd_sc_hd__o21a_1
X_13593_ _13633_/A _13634_/B VGND VGND VPWR VPWR _13593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12544_ _12544_/A VGND VGND VPWR VPWR _12544_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15332_ _15326_/Y _15330_/X _15331_/Y VGND VGND VPWR VPWR _15332_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12475_ _12465_/X _12474_/X _12465_/X _12474_/X VGND VGND VPWR VPWR _12478_/B sky130_fd_sc_hd__a2bb2o_1
X_15263_ _15218_/X _15262_/Y _15218_/X _15262_/Y VGND VGND VPWR VPWR _15264_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14214_ _14214_/A _12623_/X VGND VGND VPWR VPWR _14214_/X sky130_fd_sc_hd__or2b_1
X_11426_ _15519_/A _11429_/B VGND VGND VPWR VPWR _12586_/A sky130_fd_sc_hd__and2_1
X_15194_ _15128_/A _15128_/B _15128_/Y VGND VGND VPWR VPWR _15194_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14145_ _14145_/A VGND VGND VPWR VPWR _14145_/Y sky130_fd_sc_hd__inv_2
X_11357_ _08885_/X _11357_/B VGND VGND VPWR VPWR _11357_/X sky130_fd_sc_hd__and2b_1
XFILLER_112_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14076_ _13980_/A _13982_/X _13979_/X VGND VGND VPWR VPWR _14076_/Y sky130_fd_sc_hd__o21ai_1
X_10308_ _11759_/A _10369_/B _10307_/Y VGND VGND VPWR VPWR _10310_/A sky130_fd_sc_hd__o21ai_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13027_ _13060_/A _13025_/X _13026_/X VGND VGND VPWR VPWR _13027_/X sky130_fd_sc_hd__o21a_1
X_11288_ _12254_/A _11288_/B VGND VGND VPWR VPWR _11288_/Y sky130_fd_sc_hd__nor2_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10239_ _10239_/A _10239_/B VGND VGND VPWR VPWR _10239_/X sky130_fd_sc_hd__or2_1
XFILLER_94_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer18 rebuffer19/X VGND VGND VPWR VPWR rebuffer18/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer29 _14265_/A VGND VGND VPWR VPWR _14326_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14978_ _14971_/A _14938_/B _14938_/Y _14940_/X VGND VGND VPWR VPWR _14978_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_47_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13929_ _15400_/A _13942_/B VGND VGND VPWR VPWR _13929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09120_ _09418_/A _09123_/B VGND VGND VPWR VPWR _09120_/Y sky130_fd_sc_hd__nor2_1
X_09051_ _08712_/Y _09050_/Y _08734_/X VGND VGND VPWR VPWR _09052_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09953_ _08928_/A _09707_/Y _09627_/A _09681_/A VGND VGND VPWR VPWR _09955_/B sky130_fd_sc_hd__o22a_1
XFILLER_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _09884_/A _09884_/B VGND VGND VPWR VPWR _09885_/B sky130_fd_sc_hd__or2_1
X_08904_ _10015_/A VGND VGND VPWR VPWR _08904_/X sky130_fd_sc_hd__buf_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _09253_/B VGND VGND VPWR VPWR _10124_/A sky130_fd_sc_hd__buf_1
XFILLER_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08766_ _08765_/A _08742_/A _08765_/Y _08742_/Y VGND VGND VPWR VPWR _10132_/A sky130_fd_sc_hd__o22a_1
XFILLER_73_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08697_ _08697_/A VGND VGND VPWR VPWR _10008_/A sky130_fd_sc_hd__buf_1
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09318_ _09318_/A VGND VGND VPWR VPWR _09318_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10590_ _10590_/A VGND VGND VPWR VPWR _10590_/Y sky130_fd_sc_hd__inv_2
X_09249_ _09492_/A _09249_/B VGND VGND VPWR VPWR _10050_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12260_ _13713_/A _12259_/B _12259_/X _12166_/X VGND VGND VPWR VPWR _12260_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11211_ _11086_/X _11210_/X _11086_/X _11210_/X VGND VGND VPWR VPWR _11212_/B sky130_fd_sc_hd__a2bb2o_1
X_12191_ _13720_/A _12254_/B _12190_/Y VGND VGND VPWR VPWR _12191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11142_ _10043_/X _11142_/B VGND VGND VPWR VPWR _11142_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15950_ _15950_/A _15950_/B VGND VGND VPWR VPWR _15950_/X sky130_fd_sc_hd__or2_1
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11073_ _12135_/A _11073_/B VGND VGND VPWR VPWR _11246_/A sky130_fd_sc_hd__and2_1
XFILLER_0_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15881_ _15881_/A VGND VGND VPWR VPWR _15886_/A sky130_fd_sc_hd__inv_2
X_14901_ _14901_/A _14906_/B VGND VGND VPWR VPWR _14901_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10024_ _09250_/A _08810_/B _10073_/B _10023_/X VGND VGND VPWR VPWR _10024_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14832_ _14832_/A VGND VGND VPWR VPWR _15353_/A sky130_fd_sc_hd__buf_1
XFILLER_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14763_ _14748_/X _14762_/X _14748_/X _14762_/X VGND VGND VPWR VPWR _14833_/B sky130_fd_sc_hd__a2bb2o_1
X_11975_ _11942_/Y _11973_/X _11974_/Y VGND VGND VPWR VPWR _11975_/X sky130_fd_sc_hd__o21a_1
X_14694_ _15345_/A _14660_/B _14660_/Y VGND VGND VPWR VPWR _14694_/Y sky130_fd_sc_hd__o21ai_1
X_13714_ _12856_/A _13713_/B _13782_/A VGND VGND VPWR VPWR _13714_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10926_ _10926_/A VGND VGND VPWR VPWR _11583_/A sky130_fd_sc_hd__clkbuf_2
X_16433_ _16429_/B _16426_/A _16420_/X VGND VGND VPWR VPWR _16434_/B sky130_fd_sc_hd__a21bo_1
X_10857_ _13068_/A _10712_/B _10712_/Y VGND VGND VPWR VPWR _10857_/Y sky130_fd_sc_hd__o21ai_1
X_13645_ _13645_/A VGND VGND VPWR VPWR _13645_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16364_ _16327_/X _16363_/Y _16327_/X _16363_/Y VGND VGND VPWR VPWR _16407_/C sky130_fd_sc_hd__a2bb2o_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10788_ _11933_/A VGND VGND VPWR VPWR _13637_/A sky130_fd_sc_hd__buf_1
X_13576_ _12840_/A _13568_/B _13569_/Y _13575_/Y VGND VGND VPWR VPWR _13576_/X sky130_fd_sc_hd__o22a_1
X_16295_ _16261_/X _16294_/Y _16261_/X _16294_/Y VGND VGND VPWR VPWR _16328_/B sky130_fd_sc_hd__o2bb2a_1
X_12527_ _12633_/A _12633_/B VGND VGND VPWR VPWR _14184_/A sky130_fd_sc_hd__and2_1
X_15315_ _14580_/A _15258_/B _15258_/Y VGND VGND VPWR VPWR _15315_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15246_ _15246_/A _15246_/B VGND VGND VPWR VPWR _15246_/Y sky130_fd_sc_hd__nand2_1
X_12458_ _13883_/A _12458_/B VGND VGND VPWR VPWR _12458_/Y sky130_fd_sc_hd__nor2_1
X_11409_ _11411_/A _11409_/B VGND VGND VPWR VPWR _12320_/A sky130_fd_sc_hd__or2_1
XFILLER_125_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15177_ _15158_/X _15176_/Y _15158_/X _15176_/Y VGND VGND VPWR VPWR _15178_/B sky130_fd_sc_hd__a2bb2o_1
X_12389_ _12366_/X _12388_/Y _12366_/X _12388_/Y VGND VGND VPWR VPWR _12454_/B sky130_fd_sc_hd__a2bb2o_1
X_14128_ _14122_/X _14125_/Y _14872_/A _14127_/Y VGND VGND VPWR VPWR _14128_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14059_ _14117_/A _14057_/X _14058_/X VGND VGND VPWR VPWR _14059_/X sky130_fd_sc_hd__o21a_1
XFILLER_97_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08620_ _09457_/B VGND VGND VPWR VPWR _08717_/B sky130_fd_sc_hd__inv_2
XFILLER_94_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08551_ _08589_/A _08551_/B VGND VGND VPWR VPWR _09531_/A sky130_fd_sc_hd__or2_2
XFILLER_62_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08482_ _08276_/Y _08279_/B _08481_/Y VGND VGND VPWR VPWR _08482_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09103_ _09101_/A _08677_/B _08664_/X _09102_/Y VGND VGND VPWR VPWR _09104_/B sky130_fd_sc_hd__o22a_1
XFILLER_109_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09034_ _09551_/B _09034_/B VGND VGND VPWR VPWR _09035_/B sky130_fd_sc_hd__or2_1
XFILLER_117_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09936_ _08703_/A _09873_/A _08704_/B VGND VGND VPWR VPWR _09936_/X sky130_fd_sc_hd__o21a_1
XFILLER_100_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09867_ _08893_/X _08572_/A _09453_/Y _09866_/X VGND VGND VPWR VPWR _09867_/X sky130_fd_sc_hd__o22a_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _09251_/B VGND VGND VPWR VPWR _10126_/A sky130_fd_sc_hd__buf_1
X_09798_ _09700_/Y _09727_/A _09700_/A _09727_/Y _10940_/A VGND VGND VPWR VPWR _11907_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08749_ _08749_/A VGND VGND VPWR VPWR _08749_/Y sky130_fd_sc_hd__inv_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11760_ _10303_/A _11747_/A _10369_/B _11759_/Y VGND VGND VPWR VPWR _11761_/A sky130_fd_sc_hd__o22a_1
XFILLER_14_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10643_/A _10710_/Y _10643_/A _10710_/Y VGND VGND VPWR VPWR _10712_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11691_ _12423_/A _11691_/B VGND VGND VPWR VPWR _11691_/X sky130_fd_sc_hd__or2_1
X_13430_ _13360_/X _13429_/X _13360_/X _13429_/X VGND VGND VPWR VPWR _13430_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10642_ _10588_/Y _10640_/Y _10641_/Y VGND VGND VPWR VPWR _10643_/A sky130_fd_sc_hd__o21ai_1
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13361_ _13334_/A _13334_/B _13334_/X _13360_/X VGND VGND VPWR VPWR _13361_/X sky130_fd_sc_hd__o22a_1
X_10573_ _10671_/A _12694_/A _10572_/Y VGND VGND VPWR VPWR _10573_/X sky130_fd_sc_hd__a21o_1
X_16080_ _16027_/A _16027_/B _16027_/Y VGND VGND VPWR VPWR _16080_/X sky130_fd_sc_hd__o21a_1
X_12312_ _12312_/A _12312_/B VGND VGND VPWR VPWR _12312_/Y sky130_fd_sc_hd__nand2_1
X_13292_ _13240_/Y _13290_/Y _13291_/Y VGND VGND VPWR VPWR _13293_/A sky130_fd_sc_hd__o21ai_2
X_15100_ _15047_/X _15052_/A _15051_/X VGND VGND VPWR VPWR _15100_/X sky130_fd_sc_hd__o21a_1
Xrebuffer9 rebuffer9/A VGND VGND VPWR VPWR rebuffer9/X sky130_fd_sc_hd__dlygate4sd1_1
X_12243_ _11449_/A _12215_/B _12215_/Y _12242_/X VGND VGND VPWR VPWR _12243_/X sky130_fd_sc_hd__a2bb2o_1
X_15031_ _15079_/A _15029_/X _15030_/X VGND VGND VPWR VPWR _15031_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12174_ _12174_/A _12174_/B VGND VGND VPWR VPWR _12174_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11125_ _09919_/Y _11124_/X _09921_/A _09920_/Y _10792_/X VGND VGND VPWR VPWR _12942_/A
+ sky130_fd_sc_hd__o221a_2
X_15933_ _15956_/A _15956_/B VGND VGND VPWR VPWR _16011_/A sky130_fd_sc_hd__and2_1
X_11056_ _10908_/X _11055_/Y _10908_/X _11055_/Y VGND VGND VPWR VPWR _11076_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10007_ _08704_/B _09792_/A _09146_/X _09793_/B VGND VGND VPWR VPWR _10007_/X sky130_fd_sc_hd__a22o_1
X_15864_ _14196_/X _15846_/X _14196_/X _15846_/X VGND VGND VPWR VPWR _15898_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15795_ _15790_/Y _16227_/A _15794_/Y VGND VGND VPWR VPWR _15800_/B sky130_fd_sc_hd__o21ai_1
X_14815_ _14815_/A _14815_/B VGND VGND VPWR VPWR _14815_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14746_ _14746_/A _14746_/B VGND VGND VPWR VPWR _14746_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11958_ _11958_/A VGND VGND VPWR VPWR _13101_/A sky130_fd_sc_hd__buf_1
XFILLER_32_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10909_ _12049_/A _10909_/B VGND VGND VPWR VPWR _10909_/Y sky130_fd_sc_hd__nand2_1
X_11889_ _11889_/A _11890_/B VGND VGND VPWR VPWR _11889_/Y sky130_fd_sc_hd__nor2_1
X_14677_ _14677_/A _14677_/B VGND VGND VPWR VPWR _14677_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16416_ _16467_/Q VGND VGND VPWR VPWR _16416_/Y sky130_fd_sc_hd__inv_2
X_13628_ _13628_/A VGND VGND VPWR VPWR _13628_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16347_ _08230_/X _16469_/Q _08233_/X _16392_/B _16343_/X VGND VGND VPWR VPWR _16469_/D
+ sky130_fd_sc_hd__o221a_2
X_13559_ _13534_/X _13558_/Y _13534_/X _13558_/Y VGND VGND VPWR VPWR _13560_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16278_ _16278_/A _16277_/X VGND VGND VPWR VPWR _16278_/X sky130_fd_sc_hd__or2b_1
X_15229_ _15178_/A _15178_/B _15178_/Y _15228_/X VGND VGND VPWR VPWR _15229_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_99_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09721_ _09971_/A _09719_/Y _09720_/Y VGND VGND VPWR VPWR _09723_/B sky130_fd_sc_hd__o21ai_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09652_ _09978_/A _09652_/B VGND VGND VPWR VPWR _09652_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08603_ _09217_/A VGND VGND VPWR VPWR _10015_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09583_ _08690_/A _09017_/A _09530_/A VGND VGND VPWR VPWR _09583_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08534_ _09743_/A _08567_/B VGND VGND VPWR VPWR _08535_/A sky130_fd_sc_hd__or2_1
XFILLER_51_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08465_ _08465_/A VGND VGND VPWR VPWR _08465_/Y sky130_fd_sc_hd__inv_2
X_08396_ _09232_/A VGND VGND VPWR VPWR _08852_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09017_ _09017_/A VGND VGND VPWR VPWR _09529_/B sky130_fd_sc_hd__inv_2
XFILLER_117_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09919_ _09740_/A _09914_/Y _09861_/B VGND VGND VPWR VPWR _09919_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12930_ _12930_/A _12930_/B VGND VGND VPWR VPWR _12930_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12861_ _12792_/Y _12859_/X _12860_/Y VGND VGND VPWR VPWR _12861_/X sky130_fd_sc_hd__o21a_1
XFILLER_73_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14600_ _14600_/A _14600_/B VGND VGND VPWR VPWR _14600_/Y sky130_fd_sc_hd__nor2_1
X_11812_ _11852_/B _11811_/X _11852_/B _11811_/X VGND VGND VPWR VPWR _11848_/A sky130_fd_sc_hd__a2bb2o_1
X_15580_ _15547_/X _15579_/X _15547_/X _15579_/X VGND VGND VPWR VPWR _15581_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _13873_/A _12860_/B VGND VGND VPWR VPWR _12792_/Y sky130_fd_sc_hd__nor2_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14526_/X _14530_/X _14526_/X _14530_/X VGND VGND VPWR VPWR _14532_/B sky130_fd_sc_hd__a2bb2o_1
X_11743_ _11743_/A VGND VGND VPWR VPWR _11743_/Y sky130_fd_sc_hd__inv_2
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11671_/X _12643_/A _12642_/B VGND VGND VPWR VPWR _11674_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14454_/Y _14460_/X _14461_/Y VGND VGND VPWR VPWR _14462_/X sky130_fd_sc_hd__o21a_1
X_16201_ _16205_/A _16201_/B VGND VGND VPWR VPWR _16258_/B sky130_fd_sc_hd__or2_1
X_13413_ _14908_/A _13416_/B VGND VGND VPWR VPWR _13413_/X sky130_fd_sc_hd__and2_1
X_10625_ _11886_/A _15212_/B VGND VGND VPWR VPWR _10764_/A sky130_fd_sc_hd__or2_1
X_16132_ _16189_/A VGND VGND VPWR VPWR _16388_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14393_ _15597_/A _14391_/X _14392_/X VGND VGND VPWR VPWR _14393_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13344_ _13275_/X _13343_/Y _13275_/X _13343_/Y VGND VGND VPWR VPWR _13345_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10556_ _09421_/A _09126_/B _09126_/Y VGND VGND VPWR VPWR _10556_/X sky130_fd_sc_hd__o21a_1
X_16063_ _16052_/Y _16062_/X _16052_/Y _16062_/X VGND VGND VPWR VPWR _16121_/B sky130_fd_sc_hd__o2bb2a_1
X_13275_ _13268_/Y _13273_/X _13274_/Y VGND VGND VPWR VPWR _13275_/X sky130_fd_sc_hd__o21a_1
X_10487_ _09949_/A _10392_/B _09949_/A _10392_/B VGND VGND VPWR VPWR _10487_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12226_ _12138_/X _12225_/X _12138_/X _12225_/X VGND VGND VPWR VPWR _12227_/B sky130_fd_sc_hd__a2bb2o_1
X_15014_ _15040_/A _15040_/B VGND VGND VPWR VPWR _15064_/A sky130_fd_sc_hd__and2_1
XFILLER_123_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12157_ _12196_/A VGND VGND VPWR VPWR _13202_/A sky130_fd_sc_hd__buf_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11108_ _12196_/A VGND VGND VPWR VPWR _11276_/A sky130_fd_sc_hd__inv_2
XFILLER_96_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12088_ _12088_/A _12087_/X VGND VGND VPWR VPWR _12088_/X sky130_fd_sc_hd__or2b_1
X_15916_ _15908_/A _15908_/B _15908_/Y VGND VGND VPWR VPWR _15916_/Y sky130_fd_sc_hd__o21ai_1
X_11039_ _10912_/X _11038_/X _10912_/X _11038_/X VGND VGND VPWR VPWR _11083_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15847_ _14196_/A _15846_/X _12629_/X VGND VGND VPWR VPWR _15847_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15778_ _15778_/A _15778_/B VGND VGND VPWR VPWR _15781_/A sky130_fd_sc_hd__nor2_1
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14729_ _14729_/A _14729_/B VGND VGND VPWR VPWR _14729_/X sky130_fd_sc_hd__or2_1
X_08250_ input19/X VGND VGND VPWR VPWR _08251_/B sky130_fd_sc_hd__inv_2
XFILLER_99_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09704_ _09692_/A _09692_/B _09695_/A VGND VGND VPWR VPWR _09971_/A sky130_fd_sc_hd__a21bo_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09635_ _09635_/A VGND VGND VPWR VPWR _09635_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09566_ _09999_/A VGND VGND VPWR VPWR _09569_/A sky130_fd_sc_hd__buf_1
XFILLER_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08517_ _08516_/A _08313_/Y _08516_/Y _08313_/A VGND VGND VPWR VPWR _08518_/B sky130_fd_sc_hd__o22a_1
X_09497_ _08823_/X _09464_/X _08823_/X _09464_/X VGND VGND VPWR VPWR _09498_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_90_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08448_ _08447_/A _08318_/Y _08447_/Y _08318_/A _08441_/X VGND VGND VPWR VPWR _08543_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10410_ _09298_/A _09298_/B _09299_/A VGND VGND VPWR VPWR _10411_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08379_ _08298_/X _08378_/X _08298_/X _08378_/X VGND VGND VPWR VPWR _08662_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11390_ _08969_/X _11389_/X _08969_/X _11389_/X VGND VGND VPWR VPWR _11391_/B sky130_fd_sc_hd__a2bb2oi_2
X_10341_ _11715_/A VGND VGND VPWR VPWR _12831_/A sky130_fd_sc_hd__buf_1
XFILLER_3_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13060_ _13060_/A _13026_/X VGND VGND VPWR VPWR _13060_/X sky130_fd_sc_hd__or2b_1
X_10272_ _10272_/A VGND VGND VPWR VPWR _10272_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12011_ _13058_/A _12066_/B VGND VGND VPWR VPWR _12011_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13962_ _15420_/A _13962_/B VGND VGND VPWR VPWR _13962_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15701_ _15982_/A _14405_/B _14405_/Y VGND VGND VPWR VPWR _15701_/Y sky130_fd_sc_hd__o21ai_1
X_12913_ _10425_/A _12833_/Y _10425_/A _12833_/Y VGND VGND VPWR VPWR _12914_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13893_ _15418_/A _13960_/B VGND VGND VPWR VPWR _13893_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15632_ _15632_/A VGND VGND VPWR VPWR _15632_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12844_ _12844_/A _12844_/B VGND VGND VPWR VPWR _12844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15563_ _15563_/A _15563_/B VGND VGND VPWR VPWR _15563_/Y sky130_fd_sc_hd__nor2_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12775_ _12775_/A _12775_/B VGND VGND VPWR VPWR _12775_/Y sky130_fd_sc_hd__nand2_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _15205_/A _14514_/B VGND VGND VPWR VPWR _14514_/X sky130_fd_sc_hd__or2_1
X_11726_ _11731_/B _11725_/Y _11731_/B _11725_/Y VGND VGND VPWR VPWR _11784_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15494_ _15550_/A _15550_/B VGND VGND VPWR VPWR _15494_/X sky130_fd_sc_hd__and2_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11657_ _12788_/A _11658_/B VGND VGND VPWR VPWR _11657_/X sky130_fd_sc_hd__and2_1
X_14445_ _14467_/A _14467_/B VGND VGND VPWR VPWR _14445_/Y sky130_fd_sc_hd__nor2_1
X_14376_ _14376_/A _14376_/B VGND VGND VPWR VPWR _15661_/A sky130_fd_sc_hd__nand2_1
X_10608_ _10608_/A VGND VGND VPWR VPWR _10608_/Y sky130_fd_sc_hd__inv_2
X_11588_ _09429_/A _09750_/B _09750_/Y VGND VGND VPWR VPWR _11588_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16115_ _16067_/X _16113_/X _16155_/B VGND VGND VPWR VPWR _16119_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13327_ _13290_/A _13326_/Y _13290_/A _13326_/Y VGND VGND VPWR VPWR _13363_/B sky130_fd_sc_hd__a2bb2o_1
X_10539_ _10441_/X _10538_/B _10538_/X _10436_/X VGND VGND VPWR VPWR _10539_/X sky130_fd_sc_hd__o22a_1
X_16046_ _16046_/A _16046_/B VGND VGND VPWR VPWR _16046_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13258_ _13188_/A _13188_/B _13188_/Y VGND VGND VPWR VPWR _13258_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12209_ _14018_/A _12209_/B VGND VGND VPWR VPWR _12209_/Y sky130_fd_sc_hd__nand2_1
X_13189_ _13171_/Y _13187_/X _13188_/Y VGND VGND VPWR VPWR _13189_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09420_ _09421_/A _09421_/B VGND VGND VPWR VPWR _09420_/Y sky130_fd_sc_hd__nor2_1
X_09351_ _09351_/A VGND VGND VPWR VPWR _09351_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08302_ _08663_/B VGND VGND VPWR VPWR _08303_/A sky130_fd_sc_hd__clkbuf_2
X_09282_ _09256_/X _08963_/Y _09256_/X _08963_/Y VGND VGND VPWR VPWR _10250_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08233_ _08233_/A VGND VGND VPWR VPWR _08233_/X sky130_fd_sc_hd__buf_1
XFILLER_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08997_ _08997_/A VGND VGND VPWR VPWR _12605_/B sky130_fd_sc_hd__buf_4
XFILLER_56_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10890_ _10770_/X _10889_/Y _10770_/X _10889_/Y VGND VGND VPWR VPWR _10891_/B sky130_fd_sc_hd__a2bb2o_1
X_09618_ _09974_/A VGND VGND VPWR VPWR _09975_/A sky130_fd_sc_hd__buf_1
X_09549_ _09549_/A _09549_/B VGND VGND VPWR VPWR _09613_/B sky130_fd_sc_hd__and2_1
XFILLER_71_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12560_ _14914_/A _12344_/B _12344_/Y VGND VGND VPWR VPWR _12561_/A sky130_fd_sc_hd__o21ai_1
XFILLER_12_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12491_ _12485_/Y _12490_/Y _12485_/Y _12490_/Y VGND VGND VPWR VPWR _12494_/B sky130_fd_sc_hd__a2bb2o_1
X_11511_ _11510_/A _11510_/B _11510_/Y _10957_/X VGND VGND VPWR VPWR _11626_/A sky130_fd_sc_hd__o211a_1
XFILLER_8_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14230_ _14086_/Y _14229_/X _14086_/Y _14229_/X VGND VGND VPWR VPWR _14231_/B sky130_fd_sc_hd__a2bb2oi_1
X_11442_ _12344_/A _11446_/B VGND VGND VPWR VPWR _11442_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14161_ _14146_/X _14160_/Y _14146_/X _14160_/Y VGND VGND VPWR VPWR _14162_/B sky130_fd_sc_hd__a2bb2oi_1
X_11373_ _11391_/A _11373_/B VGND VGND VPWR VPWR _12309_/A sky130_fd_sc_hd__or2_1
XFILLER_7_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13112_ _13077_/Y _13110_/X _13111_/Y VGND VGND VPWR VPWR _13112_/X sky130_fd_sc_hd__o21a_1
X_10324_ _10324_/A VGND VGND VPWR VPWR _13528_/A sky130_fd_sc_hd__buf_1
X_14092_ _14088_/X _14090_/Y _14223_/B VGND VGND VPWR VPWR _14096_/B sky130_fd_sc_hd__o21ai_1
X_13043_ _13797_/A VGND VGND VPWR VPWR _15237_/A sky130_fd_sc_hd__buf_1
XFILLER_3_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10255_/A VGND VGND VPWR VPWR _10255_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10186_ _10244_/B _10163_/B _10163_/Y _10562_/A VGND VGND VPWR VPWR _10681_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_94_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14994_ _15765_/A VGND VGND VPWR VPWR _15752_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13945_ _13925_/Y _13943_/X _13944_/Y VGND VGND VPWR VPWR _13945_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13876_ _15110_/A _13975_/B VGND VGND VPWR VPWR _13876_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15615_ _14914_/A _15534_/B _15534_/Y VGND VGND VPWR VPWR _15617_/A sky130_fd_sc_hd__o21ai_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12827_ _12836_/A VGND VGND VPWR VPWR _15087_/A sky130_fd_sc_hd__clkbuf_2
X_15546_ _15546_/A _15546_/B VGND VGND VPWR VPWR _15586_/B sky130_fd_sc_hd__or2_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12706_/A _12706_/B _12706_/Y VGND VGND VPWR VPWR _12758_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15477_ _14806_/A _15464_/B _15464_/Y _15476_/X VGND VGND VPWR VPWR _15477_/X sky130_fd_sc_hd__a2bb2o_1
X_11709_ _12063_/A VGND VGND VPWR VPWR _13198_/A sky130_fd_sc_hd__buf_1
X_12689_ _10823_/A _12668_/A _10823_/Y _12668_/Y VGND VGND VPWR VPWR _12690_/B sky130_fd_sc_hd__o22a_1
XFILLER_30_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14428_ _11785_/X _14414_/X _11785_/X _14414_/X VGND VGND VPWR VPWR _14429_/B sky130_fd_sc_hd__a2bb2o_1
X_14359_ _13411_/Y _14358_/Y _13411_/A _14358_/A _14353_/A VGND VGND VPWR VPWR _15948_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16029_ _16027_/A _16027_/B _16027_/Y _16028_/X VGND VGND VPWR VPWR _16029_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_97_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08920_ _09541_/A _09066_/A _09235_/A _09817_/B VGND VGND VPWR VPWR _09101_/A sky130_fd_sc_hd__o22a_2
XFILLER_123_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08851_ _09677_/A VGND VGND VPWR VPWR _08916_/A sky130_fd_sc_hd__buf_1
XFILLER_111_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08782_ _08781_/A _08736_/A _08781_/Y _08736_/Y VGND VGND VPWR VPWR _10130_/A sky130_fd_sc_hd__o22a_1
XFILLER_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09403_ _09404_/A VGND VGND VPWR VPWR _09403_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09334_ _09452_/A _10130_/A VGND VGND VPWR VPWR _10044_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09265_ _09243_/X _09264_/X _09243_/X _09264_/X VGND VGND VPWR VPWR _09266_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09196_ _09198_/A VGND VGND VPWR VPWR _09196_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10040_ _10085_/A _10085_/B VGND VGND VPWR VPWR _10040_/X sky130_fd_sc_hd__and2_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11991_ _11990_/A _11990_/B _11990_/X _11925_/B VGND VGND VPWR VPWR _12080_/B sky130_fd_sc_hd__a22o_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13730_ _13730_/A _13699_/X VGND VGND VPWR VPWR _13730_/X sky130_fd_sc_hd__or2b_1
X_10942_ _12160_/A VGND VGND VPWR VPWR _13703_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15400_ _15400_/A _15400_/B VGND VGND VPWR VPWR _15400_/X sky130_fd_sc_hd__or2_1
X_10873_ _13078_/A _10729_/B _10729_/Y VGND VGND VPWR VPWR _10873_/Y sky130_fd_sc_hd__o21ai_1
X_13661_ _13699_/A _13699_/B VGND VGND VPWR VPWR _13730_/A sky130_fd_sc_hd__and2_1
X_16380_ _08230_/A _16459_/Q _08233_/A _16396_/A _16343_/A VGND VGND VPWR VPWR _16459_/D
+ sky130_fd_sc_hd__o221a_2
X_12612_ _15509_/A _12318_/B _12319_/A VGND VGND VPWR VPWR _12613_/A sky130_fd_sc_hd__o21ai_1
X_13592_ _13579_/X _13591_/Y _13579_/X _13591_/Y VGND VGND VPWR VPWR _13634_/B sky130_fd_sc_hd__a2bb2o_1
X_12543_ _12629_/A _12629_/B VGND VGND VPWR VPWR _14196_/A sky130_fd_sc_hd__and2_1
X_15331_ _15331_/A _15331_/B VGND VGND VPWR VPWR _15331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15262_ _15208_/A _15208_/B _15208_/Y VGND VGND VPWR VPWR _15262_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14213_ _14231_/A _14213_/B VGND VGND VPWR VPWR _15872_/A sky130_fd_sc_hd__or2_1
X_12474_ _12474_/A _12466_/X VGND VGND VPWR VPWR _12474_/X sky130_fd_sc_hd__or2b_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11425_ _14084_/A _11422_/B _11422_/Y _12594_/A VGND VGND VPWR VPWR _11429_/B sky130_fd_sc_hd__o2bb2a_1
X_15193_ _15193_/A _15193_/B VGND VGND VPWR VPWR _15193_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14144_ _14144_/A VGND VGND VPWR VPWR _14408_/A sky130_fd_sc_hd__inv_2
X_11356_ _12300_/A _11356_/B VGND VGND VPWR VPWR _11356_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14075_ _13997_/X _14074_/Y _13997_/X _14074_/Y VGND VGND VPWR VPWR _14075_/X sky130_fd_sc_hd__a2bb2o_1
X_10307_ _11759_/A _10369_/B VGND VGND VPWR VPWR _10307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11287_ _12360_/A VGND VGND VPWR VPWR _13042_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13026_ _14524_/A _13026_/B VGND VGND VPWR VPWR _13026_/X sky130_fd_sc_hd__or2_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10238_ _10238_/A _10238_/B VGND VGND VPWR VPWR _10238_/X sky130_fd_sc_hd__or2_1
XFILLER_121_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10169_ _10125_/A _10125_/B _10126_/B VGND VGND VPWR VPWR _10170_/B sky130_fd_sc_hd__a21bo_1
X_14977_ _14976_/Y _14954_/X _14951_/Y VGND VGND VPWR VPWR _14977_/Y sky130_fd_sc_hd__o21ai_1
X_13928_ _13841_/X _13927_/Y _13841_/X _13927_/Y VGND VGND VPWR VPWR _13942_/B sky130_fd_sc_hd__a2bb2o_1
Xrebuffer19 rebuffer20/X VGND VGND VPWR VPWR rebuffer19/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_90_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13859_ _13803_/Y _13857_/X _13858_/Y VGND VGND VPWR VPWR _13859_/X sky130_fd_sc_hd__o21a_1
X_15529_ _15529_/A _15529_/B VGND VGND VPWR VPWR _15529_/Y sky130_fd_sc_hd__nand2_1
X_09050_ _09050_/A VGND VGND VPWR VPWR _09050_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09952_ _09952_/A VGND VGND VPWR VPWR _09955_/A sky130_fd_sc_hd__inv_2
XFILLER_131_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08903_ _08684_/X _08902_/X _08684_/X _08902_/X VGND VGND VPWR VPWR _08972_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09883_/A _09883_/B VGND VGND VPWR VPWR _09884_/B sky130_fd_sc_hd__or2_1
XFILLER_112_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08834_/A VGND VGND VPWR VPWR _09253_/B sky130_fd_sc_hd__inv_2
X_08765_ _08765_/A VGND VGND VPWR VPWR _08765_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08696_ _08515_/X _08695_/Y _08515_/X _08695_/Y VGND VGND VPWR VPWR _08986_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09317_ _09263_/A _09263_/B _09263_/X _10798_/A VGND VGND VPWR VPWR _09330_/A sky130_fd_sc_hd__a22o_1
XFILLER_21_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09248_ _09248_/A VGND VGND VPWR VPWR _09263_/A sky130_fd_sc_hd__inv_2
XFILLER_119_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09179_ _09179_/A VGND VGND VPWR VPWR _09179_/Y sky130_fd_sc_hd__inv_2
X_11210_ _11210_/A _11087_/X VGND VGND VPWR VPWR _11210_/X sky130_fd_sc_hd__or2b_1
X_12190_ _12254_/A _12254_/B VGND VGND VPWR VPWR _12190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11141_ _11140_/Y _10965_/X _10976_/Y VGND VGND VPWR VPWR _11141_/X sky130_fd_sc_hd__o21a_1
X_11072_ _14430_/A _11073_/B VGND VGND VPWR VPWR _11072_/X sky130_fd_sc_hd__or2_1
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15880_ _15888_/A _15888_/B VGND VGND VPWR VPWR _15880_/Y sky130_fd_sc_hd__nor2_1
X_14900_ _14816_/X _14899_/X _14816_/X _14899_/X VGND VGND VPWR VPWR _14906_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10023_ _09456_/A _10126_/A _10069_/B _10022_/X VGND VGND VPWR VPWR _10023_/X sky130_fd_sc_hd__o22a_1
X_14831_ _14744_/X _14830_/Y _14767_/Y VGND VGND VPWR VPWR _14831_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14762_ _14762_/A _14761_/X VGND VGND VPWR VPWR _14762_/X sky130_fd_sc_hd__or2b_1
X_11974_ _13068_/A _11974_/B VGND VGND VPWR VPWR _11974_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14693_ _14739_/A _14739_/B VGND VGND VPWR VPWR _14780_/A sky130_fd_sc_hd__and2_1
XFILLER_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13713_ _13713_/A _13713_/B VGND VGND VPWR VPWR _13782_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10925_ _10925_/A VGND VGND VPWR VPWR _10925_/Y sky130_fd_sc_hd__inv_2
X_16432_ _16445_/A _16431_/Y _16445_/A _16431_/Y VGND VGND VPWR VPWR _16432_/X sky130_fd_sc_hd__a2bb2o_1
X_10856_ _12059_/A VGND VGND VPWR VPWR _10915_/A sky130_fd_sc_hd__inv_2
X_13644_ _13706_/A VGND VGND VPWR VPWR _15119_/A sky130_fd_sc_hd__buf_1
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16363_ _16328_/A _16328_/B _16328_/Y VGND VGND VPWR VPWR _16363_/Y sky130_fd_sc_hd__o21ai_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ _15339_/A _15339_/B VGND VGND VPWR VPWR _15378_/A sky130_fd_sc_hd__and2_1
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10787_ _12068_/A VGND VGND VPWR VPWR _13701_/A sky130_fd_sc_hd__buf_1
X_13575_ _13607_/A _13573_/X _13574_/X VGND VGND VPWR VPWR _13575_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16294_ _16262_/A _16328_/A _16262_/Y VGND VGND VPWR VPWR _16294_/Y sky130_fd_sc_hd__o21ai_1
X_12526_ _12525_/A _12525_/B _12525_/Y _12501_/X VGND VGND VPWR VPWR _12633_/B sky130_fd_sc_hd__o211a_1
XFILLER_75_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15245_ _15224_/X _15244_/Y _15224_/X _15244_/Y VGND VGND VPWR VPWR _15246_/B sky130_fd_sc_hd__a2bb2o_1
X_12457_ _15285_/A _12460_/B VGND VGND VPWR VPWR _12462_/A sky130_fd_sc_hd__and2_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15176_ _15110_/A _15110_/B _15110_/Y VGND VGND VPWR VPWR _15176_/Y sky130_fd_sc_hd__o21ai_1
X_11408_ _11405_/Y _11407_/Y _11405_/A _11407_/A _12605_/B VGND VGND VPWR VPWR _14084_/A
+ sky130_fd_sc_hd__o221a_4
X_14127_ _14127_/A VGND VGND VPWR VPWR _14127_/Y sky130_fd_sc_hd__inv_2
X_12388_ _13975_/A _12449_/B _12387_/Y VGND VGND VPWR VPWR _12388_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11339_ _13789_/A _11498_/B _11338_/Y VGND VGND VPWR VPWR _11339_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14058_ _14058_/A _14058_/B VGND VGND VPWR VPWR _14058_/X sky130_fd_sc_hd__or2_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13009_ _14505_/A _13008_/B _13007_/Y _13008_/Y VGND VGND VPWR VPWR _13009_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08550_ _08549_/A _08328_/Y _08549_/Y _08328_/A VGND VGND VPWR VPWR _08551_/B sky130_fd_sc_hd__o22a_1
XFILLER_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08481_ input2/X input18/X VGND VGND VPWR VPWR _08481_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09102_ _10102_/B _10098_/B VGND VGND VPWR VPWR _09102_/Y sky130_fd_sc_hd__nor2_1
X_09033_ _09549_/B _09033_/B VGND VGND VPWR VPWR _09034_/B sky130_fd_sc_hd__or2_1
XFILLER_116_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09935_ _09864_/X _09933_/X _09934_/X VGND VGND VPWR VPWR _09935_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_131_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09866_ _09454_/Y _09865_/X _09467_/X VGND VGND VPWR VPWR _09866_/X sky130_fd_sc_hd__o21a_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08817_ _08817_/A VGND VGND VPWR VPWR _09251_/B sky130_fd_sc_hd__inv_2
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09797_ _09797_/A VGND VGND VPWR VPWR _10940_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08748_ _09341_/B VGND VGND VPWR VPWR _08748_/Y sky130_fd_sc_hd__inv_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08679_/A _08679_/B VGND VGND VPWR VPWR _08679_/X sky130_fd_sc_hd__and2_1
XFILLER_26_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _13697_/A _10644_/B _10644_/Y VGND VGND VPWR VPWR _10710_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11690_ _12423_/B VGND VGND VPWR VPWR _11691_/B sky130_fd_sc_hd__inv_2
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10641_ _11904_/A _10641_/B VGND VGND VPWR VPWR _10641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13360_ _13337_/A _13337_/B _13337_/X _13359_/X VGND VGND VPWR VPWR _13360_/X sky130_fd_sc_hd__o22a_1
X_10572_ _10671_/A _11918_/A VGND VGND VPWR VPWR _10572_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12311_ _12243_/X _12310_/Y _12243_/X _12310_/Y VGND VGND VPWR VPWR _12312_/B sky130_fd_sc_hd__a2bb2o_1
X_13291_ _14735_/A _13291_/B VGND VGND VPWR VPWR _13291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12242_ _12218_/A _12218_/B _12218_/Y _12241_/X VGND VGND VPWR VPWR _12242_/X sky130_fd_sc_hd__a2bb2o_1
X_15030_ _15030_/A _15030_/B VGND VGND VPWR VPWR _15030_/X sky130_fd_sc_hd__or2_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12173_ _12172_/A _12172_/B _12172_/X _12087_/B VGND VGND VPWR VPWR _12266_/B sky130_fd_sc_hd__a22o_1
XFILLER_96_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11124_ _09918_/A _09918_/B _09921_/A VGND VGND VPWR VPWR _11124_/X sky130_fd_sc_hd__o21ba_1
X_15932_ _15893_/X _15931_/Y _15893_/X _15931_/Y VGND VGND VPWR VPWR _15956_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11055_ _12049_/A _10909_/B _10909_/Y VGND VGND VPWR VPWR _11055_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10006_ _11710_/A VGND VGND VPWR VPWR _13525_/A sky130_fd_sc_hd__buf_1
X_15863_ _15863_/A VGND VGND VPWR VPWR _15898_/A sky130_fd_sc_hd__inv_2
XFILLER_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15794_ _16094_/A _15794_/B VGND VGND VPWR VPWR _15794_/Y sky130_fd_sc_hd__nand2_1
X_14814_ _13937_/X _14813_/Y _13937_/X _14813_/Y VGND VGND VPWR VPWR _14815_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14745_ _14745_/A VGND VGND VPWR VPWR _15351_/A sky130_fd_sc_hd__buf_1
X_11957_ _11964_/A _11964_/B VGND VGND VPWR VPWR _12038_/A sky130_fd_sc_hd__and2_1
X_10908_ _13833_/A _10907_/B _11065_/A _10907_/Y VGND VGND VPWR VPWR _10908_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16415_ _16415_/A VGND VGND VPWR VPWR _16415_/X sky130_fd_sc_hd__buf_1
X_11888_ _10623_/A _11887_/X _10623_/A _11887_/X VGND VGND VPWR VPWR _11890_/B sky130_fd_sc_hd__a2bb2o_1
X_14676_ _14671_/X _14675_/X _14671_/X _14675_/X VGND VGND VPWR VPWR _14677_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13627_ _13599_/Y _13624_/Y _13626_/Y VGND VGND VPWR VPWR _13628_/A sky130_fd_sc_hd__o21ai_2
X_10839_ _12068_/A _10935_/B VGND VGND VPWR VPWR _10839_/Y sky130_fd_sc_hd__nand2_1
X_16346_ _16337_/X _16345_/Y _16337_/X _16345_/Y VGND VGND VPWR VPWR _16392_/B sky130_fd_sc_hd__a2bb2o_1
X_13558_ _15034_/A _13522_/B _13522_/Y VGND VGND VPWR VPWR _13558_/Y sky130_fd_sc_hd__o21ai_1
X_16277_ _16277_/A _16277_/B VGND VGND VPWR VPWR _16277_/X sky130_fd_sc_hd__or2_1
X_12509_ _12509_/A _12509_/B VGND VGND VPWR VPWR _12509_/Y sky130_fd_sc_hd__nand2_1
X_15228_ _15181_/A _15181_/B _15181_/Y _15227_/X VGND VGND VPWR VPWR _15228_/X sky130_fd_sc_hd__a2bb2o_1
X_13489_ _10960_/Y _11997_/A _10829_/Y _13488_/X VGND VGND VPWR VPWR _13489_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15159_ _15110_/A _15110_/B _15110_/Y _15158_/X VGND VGND VPWR VPWR _15159_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_101_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09720_ _09720_/A _09720_/B VGND VGND VPWR VPWR _09720_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09651_ _09647_/Y _10722_/A _09650_/Y VGND VGND VPWR VPWR _09651_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08602_ _09456_/B VGND VGND VPWR VPWR _09549_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09582_ _09992_/A VGND VGND VPWR VPWR _09993_/A sky130_fd_sc_hd__buf_1
XFILLER_82_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08533_ _09861_/A VGND VGND VPWR VPWR _09743_/A sky130_fd_sc_hd__inv_2
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08464_ _08464_/A VGND VGND VPWR VPWR _08464_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08395_ _08934_/A VGND VGND VPWR VPWR _09232_/A sky130_fd_sc_hd__inv_2
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09016_ _08770_/A _09015_/X _09015_/X _08546_/Y VGND VGND VPWR VPWR _09017_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09918_ _09918_/A _09918_/B VGND VGND VPWR VPWR _09921_/A sky130_fd_sc_hd__and2_1
XFILLER_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09849_ _09693_/A _09844_/Y _09803_/B VGND VGND VPWR VPWR _09849_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12860_ _13873_/A _12860_/B VGND VGND VPWR VPWR _12860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11811_/A _11810_/X VGND VGND VPWR VPWR _11811_/X sky130_fd_sc_hd__or2b_1
XFILLER_27_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14529_/A _14529_/B _14529_/Y VGND VGND VPWR VPWR _14530_/X sky130_fd_sc_hd__a21o_1
X_12791_ _12784_/X _12790_/Y _12784_/X _12790_/Y VGND VGND VPWR VPWR _12860_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11742_/A _11742_/B VGND VGND VPWR VPWR _11742_/X sky130_fd_sc_hd__or2_1
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _15554_/A _11673_/B VGND VGND VPWR VPWR _12642_/B sky130_fd_sc_hd__or2_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14461_/A _14461_/B VGND VGND VPWR VPWR _14461_/Y sky130_fd_sc_hd__nand2_1
X_16200_ _16103_/X _16199_/X _16103_/X _16199_/X VGND VGND VPWR VPWR _16201_/B sky130_fd_sc_hd__o2bb2a_1
X_14392_ _15962_/A _14392_/B VGND VGND VPWR VPWR _14392_/X sky130_fd_sc_hd__or2_1
X_13412_ _14901_/A _13408_/B _13408_/X _13411_/Y VGND VGND VPWR VPWR _13416_/B sky130_fd_sc_hd__o22a_1
X_10624_ _12041_/A VGND VGND VPWR VPWR _15212_/B sky130_fd_sc_hd__inv_2
X_16131_ _16205_/A VGND VGND VPWR VPWR _16189_/A sky130_fd_sc_hd__buf_1
X_13343_ _14725_/A _13276_/B _13276_/Y VGND VGND VPWR VPWR _13343_/Y sky130_fd_sc_hd__o21ai_1
X_10555_ _10554_/Y _10454_/X _10465_/Y VGND VGND VPWR VPWR _10555_/X sky130_fd_sc_hd__o21a_1
X_16062_ _15998_/X _16062_/B VGND VGND VPWR VPWR _16062_/X sky130_fd_sc_hd__and2b_1
X_13274_ _13274_/A _13274_/B VGND VGND VPWR VPWR _13274_/Y sky130_fd_sc_hd__nand2_1
X_10486_ _11841_/A VGND VGND VPWR VPWR _13625_/A sky130_fd_sc_hd__buf_1
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12225_ _12225_/A _12139_/X VGND VGND VPWR VPWR _12225_/X sky130_fd_sc_hd__or2b_1
X_15013_ _11926_/X _15003_/X _11926_/X _15003_/X VGND VGND VPWR VPWR _15040_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12156_ _12155_/Y _12064_/X _12104_/Y VGND VGND VPWR VPWR _12156_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11107_ _11106_/A _11105_/Y _11106_/Y _11105_/A _11583_/A VGND VGND VPWR VPWR _12196_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_77_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12087_ _12087_/A _12087_/B VGND VGND VPWR VPWR _12087_/X sky130_fd_sc_hd__or2_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15915_ _15972_/A _15972_/B VGND VGND VPWR VPWR _15993_/A sky130_fd_sc_hd__and2_1
XFILLER_110_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11038_ _10875_/A _10875_/B _10875_/A _10875_/B VGND VGND VPWR VPWR _11038_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15846_ _14202_/A _15845_/X _12627_/X VGND VGND VPWR VPWR _15846_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15777_ _15782_/A _15782_/B VGND VGND VPWR VPWR _16245_/A sky130_fd_sc_hd__and2_1
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12989_ _14489_/A _13018_/B VGND VGND VPWR VPWR _13080_/A sky130_fd_sc_hd__and2_1
XFILLER_52_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14728_ _14804_/A _14726_/Y _14727_/X VGND VGND VPWR VPWR _14728_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14659_ _14618_/Y _14657_/X _14658_/Y VGND VGND VPWR VPWR _14659_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16329_ _16296_/Y _16327_/X _16328_/Y VGND VGND VPWR VPWR _16329_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09703_ _09703_/A VGND VGND VPWR VPWR _09723_/A sky130_fd_sc_hd__inv_2
XFILLER_114_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09634_ _09629_/B _09633_/Y _09629_/B _09633_/Y VGND VGND VPWR VPWR _09635_/A sky130_fd_sc_hd__a2bb2o_1
X_09565_ _09563_/Y _09564_/X _09563_/Y _09564_/X VGND VGND VPWR VPWR _09999_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08516_ _08516_/A VGND VGND VPWR VPWR _08516_/Y sky130_fd_sc_hd__inv_2
X_09496_ _09496_/A _09496_/B VGND VGND VPWR VPWR _09496_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08447_ _08447_/A VGND VGND VPWR VPWR _08447_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08378_ input7/X _08235_/B _08238_/B _08465_/A VGND VGND VPWR VPWR _08378_/X sky130_fd_sc_hd__o22a_2
XFILLER_99_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10340_ _08929_/B _10339_/Y _08928_/A _10277_/Y _10446_/A VGND VGND VPWR VPWR _11715_/A
+ sky130_fd_sc_hd__o221a_1
X_10271_ _09298_/A _10230_/B _10231_/A VGND VGND VPWR VPWR _10272_/A sky130_fd_sc_hd__o21ai_1
X_12010_ _12069_/A _12009_/Y _12069_/A _12009_/Y VGND VGND VPWR VPWR _12066_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13961_ _13893_/Y _13959_/X _13960_/Y VGND VGND VPWR VPWR _13961_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15700_ _15700_/A _15700_/B VGND VGND VPWR VPWR _15991_/A sky130_fd_sc_hd__or2_1
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12912_ _13610_/A VGND VGND VPWR VPWR _13003_/A sky130_fd_sc_hd__buf_1
XFILLER_59_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13892_ _13859_/X _13891_/Y _13859_/X _13891_/Y VGND VGND VPWR VPWR _13960_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15631_ _14910_/A _15524_/B _15524_/Y VGND VGND VPWR VPWR _15633_/A sky130_fd_sc_hd__o21ai_1
XFILLER_104_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12843_ _12819_/Y _12841_/X _12842_/Y VGND VGND VPWR VPWR _12843_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15562_ _15559_/X _15561_/X _15559_/X _15561_/X VGND VGND VPWR VPWR _15562_/X sky130_fd_sc_hd__a2bb2o_1
X_12774_ _12744_/Y _12772_/X _12773_/Y VGND VGND VPWR VPWR _12774_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15493_ _15484_/X _15492_/X _15484_/X _15492_/X VGND VGND VPWR VPWR _15550_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14561_/A _14511_/X _14512_/X VGND VGND VPWR VPWR _14513_/X sky130_fd_sc_hd__o21a_1
X_11725_ _11724_/A _11730_/A _11724_/Y VGND VGND VPWR VPWR _11725_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _14435_/X _14443_/X _14435_/X _14443_/X VGND VGND VPWR VPWR _14467_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11656_ _11580_/X _11655_/X _11580_/X _11655_/X VGND VGND VPWR VPWR _11658_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14375_ _14375_/A VGND VGND VPWR VPWR _14375_/Y sky130_fd_sc_hd__inv_2
X_11587_ _11587_/A _11587_/B VGND VGND VPWR VPWR _12443_/A sky130_fd_sc_hd__or2_2
X_10607_ _09407_/A _09709_/B _09709_/Y VGND VGND VPWR VPWR _10608_/A sky130_fd_sc_hd__o21ai_1
XFILLER_128_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16114_ _16114_/A _16114_/B VGND VGND VPWR VPWR _16155_/B sky130_fd_sc_hd__or2_1
X_13326_ _14735_/A _13291_/B _13291_/Y VGND VGND VPWR VPWR _13326_/Y sky130_fd_sc_hd__o21ai_1
X_10538_ _11028_/A _10538_/B VGND VGND VPWR VPWR _10538_/X sky130_fd_sc_hd__and2_1
X_16045_ _16004_/Y _16043_/X _16044_/Y VGND VGND VPWR VPWR _16045_/X sky130_fd_sc_hd__o21a_1
X_13257_ _14425_/A VGND VGND VPWR VPWR _14727_/A sky130_fd_sc_hd__buf_1
XFILLER_89_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12208_ _12150_/X _12207_/X _12150_/X _12207_/X VGND VGND VPWR VPWR _12209_/B sky130_fd_sc_hd__a2bb2o_1
X_10469_ _10469_/A VGND VGND VPWR VPWR _10469_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13188_ _13188_/A _13188_/B VGND VGND VPWR VPWR _13188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12139_ _14427_/A _12139_/B VGND VGND VPWR VPWR _12139_/X sky130_fd_sc_hd__or2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15829_ _15824_/X _15828_/Y _15824_/X _15828_/Y VGND VGND VPWR VPWR _15829_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09350_ _09527_/A _09743_/A VGND VGND VPWR VPWR _09351_/A sky130_fd_sc_hd__or2_1
XFILLER_33_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09281_ _09240_/Y _09280_/X _09240_/Y _09280_/X VGND VGND VPWR VPWR _09946_/A sky130_fd_sc_hd__a2bb2o_2
X_08301_ _08400_/B VGND VGND VPWR VPWR _08663_/B sky130_fd_sc_hd__inv_2
X_08232_ _08232_/A VGND VGND VPWR VPWR _08233_/A sky130_fd_sc_hd__buf_1
XFILLER_119_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08996_ _08988_/X _08995_/X _08988_/X _08995_/X VGND VGND VPWR VPWR _08997_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09617_ _09508_/X _09616_/X _09508_/X _09616_/X VGND VGND VPWR VPWR _09974_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09548_ _09648_/A _09546_/Y _09648_/B VGND VGND VPWR VPWR _09548_/X sky130_fd_sc_hd__o21ba_1
X_11510_ _11510_/A _11510_/B VGND VGND VPWR VPWR _11510_/Y sky130_fd_sc_hd__nand2_1
X_09479_ _09448_/Y _09477_/X _09478_/X VGND VGND VPWR VPWR _09520_/S sky130_fd_sc_hd__o21ai_1
X_12490_ _12486_/A _12486_/B _12486_/Y VGND VGND VPWR VPWR _12490_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11441_ _11436_/Y _12564_/A _11440_/Y VGND VGND VPWR VPWR _11446_/B sky130_fd_sc_hd__o21ai_2
XFILLER_125_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14160_ _13450_/A _14149_/B _14149_/Y VGND VGND VPWR VPWR _14160_/Y sky130_fd_sc_hd__a21oi_1
X_11372_ _08975_/X _11371_/X _08975_/X _11371_/X VGND VGND VPWR VPWR _11373_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_125_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13111_ _15255_/A _13111_/B VGND VGND VPWR VPWR _13111_/Y sky130_fd_sc_hd__nand2_1
X_10323_ _11776_/A VGND VGND VPWR VPWR _10324_/A sky130_fd_sc_hd__inv_2
XFILLER_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14091_ _14091_/A _14091_/B VGND VGND VPWR VPWR _14223_/B sky130_fd_sc_hd__or2_1
XFILLER_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13042_ _13042_/A VGND VGND VPWR VPWR _13797_/A sky130_fd_sc_hd__inv_2
X_10254_ _10254_/A _10254_/B VGND VGND VPWR VPWR _10255_/A sky130_fd_sc_hd__nand2_1
X_10185_ _10469_/A _10167_/B _10167_/Y _10462_/A VGND VGND VPWR VPWR _10562_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14993_ _15778_/B VGND VGND VPWR VPWR _15765_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13944_ _15402_/A _13944_/B VGND VGND VPWR VPWR _13944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13875_ _13869_/X _13874_/X _13869_/X _13874_/X VGND VGND VPWR VPWR _13975_/B sky130_fd_sc_hd__a2bb2o_1
X_15614_ _15677_/A _15677_/B VGND VGND VPWR VPWR _15614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12826_ _12826_/A VGND VGND VPWR VPWR _12836_/A sky130_fd_sc_hd__inv_2
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15545_ _15503_/X _15543_/X _15593_/B VGND VGND VPWR VPWR _15545_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _15028_/A VGND VGND VPWR VPWR _12763_/A sky130_fd_sc_hd__inv_2
X_11708_ _11566_/A _11566_/B _11566_/Y _11707_/X VGND VGND VPWR VPWR _12639_/A sky130_fd_sc_hd__o211a_1
X_15476_ _15467_/A _15467_/B _15467_/Y _15475_/X VGND VGND VPWR VPWR _15476_/X sky130_fd_sc_hd__a2bb2o_1
X_12688_ _12688_/A _12688_/B VGND VGND VPWR VPWR _12688_/Y sky130_fd_sc_hd__nor2_1
X_14427_ _14427_/A _14427_/B VGND VGND VPWR VPWR _14427_/X sky130_fd_sc_hd__and2_1
X_11639_ _11638_/Y _11499_/X _11543_/Y VGND VGND VPWR VPWR _11639_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14358_ _14358_/A VGND VGND VPWR VPWR _14358_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13309_ _14068_/A _13309_/B VGND VGND VPWR VPWR _13309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14289_ _14295_/A _14287_/X _14288_/X VGND VGND VPWR VPWR _14289_/X sky130_fd_sc_hd__o21a_1
X_16028_ _16028_/A _16028_/B VGND VGND VPWR VPWR _16028_/X sky130_fd_sc_hd__or2_1
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08850_ _08852_/A VGND VGND VPWR VPWR _09503_/A sky130_fd_sc_hd__buf_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08781_ _08781_/A VGND VGND VPWR VPWR _08781_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09402_ _09817_/B _09707_/B _09401_/Y VGND VGND VPWR VPWR _09404_/A sky130_fd_sc_hd__a21oi_1
XFILLER_80_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09333_ _09333_/A _10131_/A VGND VGND VPWR VPWR _10041_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09264_ _09467_/B _09857_/A _09212_/A VGND VGND VPWR VPWR _09264_/X sky130_fd_sc_hd__o21a_1
X_09195_ _09167_/Y _09194_/Y _09167_/Y _09194_/Y VGND VGND VPWR VPWR _09198_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08979_ _08890_/X _08977_/X _11364_/B VGND VGND VPWR VPWR _08979_/X sky130_fd_sc_hd__o21a_1
X_11990_ _11990_/A _11990_/B VGND VGND VPWR VPWR _11990_/X sky130_fd_sc_hd__or2_1
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10941_ _09967_/Y _10939_/A _10081_/A _10939_/Y _11590_/A VGND VGND VPWR VPWR _12160_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13660_ _13636_/A _13659_/Y _13636_/A _13659_/Y VGND VGND VPWR VPWR _13699_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12611_ _14082_/A VGND VGND VPWR VPWR _15509_/A sky130_fd_sc_hd__buf_1
X_10872_ _10875_/A VGND VGND VPWR VPWR _14627_/A sky130_fd_sc_hd__buf_1
XFILLER_44_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13591_ _13552_/A _13552_/B _13553_/A VGND VGND VPWR VPWR _13591_/Y sky130_fd_sc_hd__o21ai_1
X_12542_ _12541_/A _12541_/B _12541_/Y _12501_/A VGND VGND VPWR VPWR _12629_/B sky130_fd_sc_hd__o211a_1
X_15330_ _15329_/A _15329_/B _12043_/Y _15329_/Y VGND VGND VPWR VPWR _15330_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_12_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15261_ _15261_/A _15261_/B VGND VGND VPWR VPWR _15261_/Y sky130_fd_sc_hd__nand2_1
X_12473_ _12431_/X _12472_/X _12431_/X _12472_/X VGND VGND VPWR VPWR _12473_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_12_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14212_ _14100_/Y _14211_/X _14100_/Y _14211_/X VGND VGND VPWR VPWR _14213_/B sky130_fd_sc_hd__a2bb2oi_1
X_11424_ _11251_/X _11423_/Y _11251_/X _11423_/Y VGND VGND VPWR VPWR _12594_/A sky130_fd_sc_hd__a2bb2o_1
X_15192_ _15153_/X _15191_/Y _15153_/X _15191_/Y VGND VGND VPWR VPWR _15193_/B sky130_fd_sc_hd__a2bb2o_1
X_14143_ _14144_/A _14145_/A VGND VGND VPWR VPWR _14143_/Y sky130_fd_sc_hd__nor2_1
X_11355_ _11261_/X _11354_/Y _11261_/X _11354_/Y VGND VGND VPWR VPWR _11356_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14074_ _13999_/X _14073_/X _13999_/X _14073_/X VGND VGND VPWR VPWR _14074_/Y sky130_fd_sc_hd__a2bb2oi_1
X_11286_ _11587_/A _11286_/B VGND VGND VPWR VPWR _12360_/A sky130_fd_sc_hd__or2_1
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10306_ _10182_/A _10305_/A _10182_/Y _10305_/Y _10463_/A VGND VGND VPWR VPWR _10369_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13025_ _13065_/A _13023_/X _13024_/X VGND VGND VPWR VPWR _13025_/X sky130_fd_sc_hd__o21a_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ _11574_/A _10237_/B VGND VGND VPWR VPWR _10237_/X sky130_fd_sc_hd__or2_1
XFILLER_121_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10168_ _10112_/A _10112_/B _10113_/A VGND VGND VPWR VPWR _10251_/A sky130_fd_sc_hd__a21bo_1
XFILLER_86_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14976_ _14976_/A _14976_/B VGND VGND VPWR VPWR _14976_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10099_ _10099_/A _10099_/B VGND VGND VPWR VPWR _10110_/A sky130_fd_sc_hd__or2_1
X_13927_ _14635_/A _13842_/B _13842_/Y VGND VGND VPWR VPWR _13927_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13858_ _14664_/A _13858_/B VGND VGND VPWR VPWR _13858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13789_ _13789_/A _13865_/B VGND VGND VPWR VPWR _13789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12809_ _12772_/X _12808_/Y _12772_/X _12808_/Y VGND VGND VPWR VPWR _12848_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15528_ _15477_/X _15527_/Y _15477_/X _15527_/Y VGND VGND VPWR VPWR _15624_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15459_ _15459_/A _15404_/X VGND VGND VPWR VPWR _15459_/X sky130_fd_sc_hd__or2b_1
XFILLER_30_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09951_ _10216_/A VGND VGND VPWR VPWR _09951_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08902_ _09551_/A _08596_/A _08598_/A VGND VGND VPWR VPWR _08902_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _09882_/A _09882_/B VGND VGND VPWR VPWR _09883_/B sky130_fd_sc_hd__or2_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _09228_/A VGND VGND VPWR VPWR _10018_/A sky130_fd_sc_hd__buf_1
XFILLER_111_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _09331_/A _09476_/B _08709_/Y VGND VGND VPWR VPWR _08765_/A sky130_fd_sc_hd__a21oi_2
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08695_ _08871_/A _08693_/X _08871_/B VGND VGND VPWR VPWR _08695_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09316_ _09269_/A _09269_/B _09269_/X _10660_/A VGND VGND VPWR VPWR _10798_/A sky130_fd_sc_hd__a22o_1
X_09247_ _09244_/X _09246_/X _09244_/X _09246_/X VGND VGND VPWR VPWR _09248_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09178_ _09527_/B _09155_/B _09156_/B VGND VGND VPWR VPWR _09179_/A sky130_fd_sc_hd__a21bo_1
Xoutput34 _16472_/Q VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__clkbuf_2
X_11140_ _12174_/A _11140_/B VGND VGND VPWR VPWR _11140_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11071_ _11065_/A _11070_/X _11065_/A _11070_/X VGND VGND VPWR VPWR _11073_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10022_ _09252_/A _10125_/A _10065_/B _10021_/X VGND VGND VPWR VPWR _10022_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14830_ _15351_/A _14830_/B VGND VGND VPWR VPWR _14830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11973_ _11945_/Y _11971_/X _11972_/Y VGND VGND VPWR VPWR _11973_/X sky130_fd_sc_hd__o21a_1
X_14761_ _15181_/A _14761_/B VGND VGND VPWR VPWR _14761_/X sky130_fd_sc_hd__or2_1
XFILLER_56_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14692_ _14661_/X _14691_/Y _14661_/X _14691_/Y VGND VGND VPWR VPWR _14739_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13712_ _13540_/X _13711_/Y _13540_/X _13711_/Y VGND VGND VPWR VPWR _13713_/B sky130_fd_sc_hd__a2bb2o_1
X_10924_ _09436_/A _09436_/B _09436_/Y VGND VGND VPWR VPWR _10925_/A sky130_fd_sc_hd__o21ai_1
X_16431_ _16437_/D _16419_/B _16445_/B VGND VGND VPWR VPWR _16431_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13643_ _13587_/Y _13640_/Y _13642_/Y VGND VGND VPWR VPWR _13705_/A sky130_fd_sc_hd__o21ai_2
X_10855_ _09272_/A _10854_/A _09275_/A _10854_/Y _10926_/A VGND VGND VPWR VPWR _12059_/A
+ sky130_fd_sc_hd__a221o_2
X_16362_ _16357_/X _16465_/Q _16358_/X _16407_/D _16361_/X VGND VGND VPWR VPWR _16465_/D
+ sky130_fd_sc_hd__o221a_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13574_ _14429_/A _13574_/B VGND VGND VPWR VPWR _13574_/X sky130_fd_sc_hd__or2_1
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12525_ _12525_/A _12525_/B VGND VGND VPWR VPWR _12525_/Y sky130_fd_sc_hd__nand2_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15313_ _15276_/X _15312_/Y _15276_/X _15312_/Y VGND VGND VPWR VPWR _15339_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10786_ _09968_/Y _10785_/A _10079_/A _10785_/Y _10940_/A VGND VGND VPWR VPWR _12068_/A
+ sky130_fd_sc_hd__a221o_2
X_16293_ _16330_/A _16330_/B VGND VGND VPWR VPWR _16293_/Y sky130_fd_sc_hd__nor2_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15244_ _15190_/A _15190_/B _15190_/Y VGND VGND VPWR VPWR _15244_/Y sky130_fd_sc_hd__o21ai_1
X_12456_ _12453_/X _12480_/A _12453_/X _12480_/A VGND VGND VPWR VPWR _12460_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15175_ _15556_/A _15556_/B _15174_/Y VGND VGND VPWR VPWR _15175_/Y sky130_fd_sc_hd__o21ai_1
X_12387_ _12387_/A _12449_/B VGND VGND VPWR VPWR _12387_/Y sky130_fd_sc_hd__nand2_1
X_11407_ _11407_/A VGND VGND VPWR VPWR _11407_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14126_ _14126_/A VGND VGND VPWR VPWR _14872_/A sky130_fd_sc_hd__inv_2
X_11338_ _12365_/A _11498_/B VGND VGND VPWR VPWR _11338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14057_ _14077_/A _14055_/X _14056_/X VGND VGND VPWR VPWR _14057_/X sky130_fd_sc_hd__o21a_1
X_11269_ _11269_/A _11269_/B VGND VGND VPWR VPWR _11269_/Y sky130_fd_sc_hd__nand2_1
X_13008_ _14505_/A _13008_/B VGND VGND VPWR VPWR _13008_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14959_ _14831_/X _14958_/Y _14854_/Y VGND VGND VPWR VPWR _14959_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08480_ input26/X input10/X VGND VGND VPWR VPWR _08480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09101_ _09101_/A VGND VGND VPWR VPWR _10102_/B sky130_fd_sc_hd__inv_2
X_09032_ _09547_/B _09032_/B VGND VGND VPWR VPWR _09033_/B sky130_fd_sc_hd__or2_1
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09934_ _09863_/X _09932_/X _09863_/X _09932_/X VGND VGND VPWR VPWR _09934_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09865_ _08904_/X _08597_/A _09455_/Y _09812_/X VGND VGND VPWR VPWR _09865_/X sky130_fd_sc_hd__o22a_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08816_ _10016_/A VGND VGND VPWR VPWR _08819_/A sky130_fd_sc_hd__buf_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09796_ _10618_/A VGND VGND VPWR VPWR _09797_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08747_ _08708_/Y _08745_/Y _08746_/X VGND VGND VPWR VPWR _09341_/B sky130_fd_sc_hd__o21ai_2
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08678_/A VGND VGND VPWR VPWR _08678_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10640_/A VGND VGND VPWR VPWR _10640_/Y sky130_fd_sc_hd__inv_2
X_10571_ _11918_/A VGND VGND VPWR VPWR _12694_/A sky130_fd_sc_hd__buf_1
X_12310_ _14021_/A _12212_/B _12212_/Y VGND VGND VPWR VPWR _12310_/Y sky130_fd_sc_hd__o21ai_1
X_13290_ _13290_/A VGND VGND VPWR VPWR _13290_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12241_ _12221_/A _12221_/B _12221_/Y _12240_/X VGND VGND VPWR VPWR _12241_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12172_ _12172_/A _12172_/B VGND VGND VPWR VPWR _12172_/X sky130_fd_sc_hd__or2_1
XFILLER_122_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11123_ _11122_/Y _10945_/X _10992_/Y VGND VGND VPWR VPWR _11123_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15931_ _15894_/A _15894_/B _15894_/Y VGND VGND VPWR VPWR _15931_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11054_ _15084_/A VGND VGND VPWR VPWR _12137_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10005_ _09963_/A _09962_/Y _09963_/Y _09962_/A _10446_/A VGND VGND VPWR VPWR _11710_/A
+ sky130_fd_sc_hd__o221a_1
X_15862_ _15900_/A _15900_/B VGND VGND VPWR VPWR _15862_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15793_ _15793_/A VGND VGND VPWR VPWR _16094_/A sky130_fd_sc_hd__buf_1
XFILLER_123_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14813_ _14722_/A _14722_/B _14722_/Y VGND VGND VPWR VPWR _14813_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14744_ _14663_/X _14743_/Y _14687_/Y VGND VGND VPWR VPWR _14744_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11956_ _11891_/X _11955_/Y _11891_/X _11955_/Y VGND VGND VPWR VPWR _11964_/B sky130_fd_sc_hd__a2bb2o_1
X_10907_ _12047_/A _10907_/B VGND VGND VPWR VPWR _10907_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16414_ _16437_/D _16473_/Q VGND VGND VPWR VPWR _16415_/A sky130_fd_sc_hd__or2_1
X_11887_ _13610_/A _11833_/B _11833_/Y VGND VGND VPWR VPWR _11887_/X sky130_fd_sc_hd__a21o_1
X_14675_ _14674_/A _14674_/B _14674_/Y VGND VGND VPWR VPWR _14675_/X sky130_fd_sc_hd__a21o_1
X_13626_ _15134_/A _13626_/B VGND VGND VPWR VPWR _13626_/Y sky130_fd_sc_hd__nand2_1
X_10838_ _10790_/X _10837_/Y _10790_/X _10837_/Y VGND VGND VPWR VPWR _10935_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16345_ _16338_/A _16338_/B _16338_/Y VGND VGND VPWR VPWR _16345_/Y sky130_fd_sc_hd__o21ai_1
X_10769_ _14564_/A _10769_/B VGND VGND VPWR VPWR _10769_/X sky130_fd_sc_hd__or2_1
X_13557_ _13557_/A VGND VGND VPWR VPWR _13557_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16276_ _16277_/A _16277_/B VGND VGND VPWR VPWR _16278_/A sky130_fd_sc_hd__and2_1
X_12508_ _13446_/A _12300_/B _12300_/Y VGND VGND VPWR VPWR _12509_/B sky130_fd_sc_hd__o21a_1
X_13488_ _10807_/Y _11925_/A _10691_/Y _13487_/X VGND VGND VPWR VPWR _13488_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15227_ _15184_/A _15184_/B _15184_/Y _15226_/X VGND VGND VPWR VPWR _15227_/X sky130_fd_sc_hd__a2bb2o_1
X_12439_ _13463_/A _12439_/B VGND VGND VPWR VPWR _12439_/X sky130_fd_sc_hd__and2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15158_ _15113_/A _15113_/B _15113_/Y _15157_/X VGND VGND VPWR VPWR _15158_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14109_ _14109_/A VGND VGND VPWR VPWR _15455_/A sky130_fd_sc_hd__buf_1
X_15089_ _12137_/A _15084_/B _15084_/Y _15088_/X VGND VGND VPWR VPWR _15089_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09650_ _09975_/A _09650_/B VGND VGND VPWR VPWR _09650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08601_ _08650_/A _08601_/B VGND VGND VPWR VPWR _09456_/B sky130_fd_sc_hd__or2_1
XFILLER_94_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09581_ _09514_/X _09580_/X _09514_/X _09580_/X VGND VGND VPWR VPWR _09992_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08532_ _08532_/A _08532_/B VGND VGND VPWR VPWR _09861_/A sky130_fd_sc_hd__or2_2
XFILLER_63_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08463_ _08521_/B _08459_/Y _09448_/A VGND VGND VPWR VPWR _08464_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08394_ _08662_/A _08394_/B VGND VGND VPWR VPWR _08934_/A sky130_fd_sc_hd__or2_2
XFILLER_50_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09015_ _08778_/A _09014_/Y _08555_/B VGND VGND VPWR VPWR _09015_/X sky130_fd_sc_hd__o21ba_1
XFILLER_105_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09917_ _10947_/B _09916_/X VGND VGND VPWR VPWR _09918_/B sky130_fd_sc_hd__or2b_1
XFILLER_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09848_ _09848_/A _09848_/B VGND VGND VPWR VPWR _09851_/A sky130_fd_sc_hd__and2_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09779_ _09779_/A _09779_/B VGND VGND VPWR VPWR _09779_/Y sky130_fd_sc_hd__nand2_1
X_12790_ _12785_/A _12785_/B _12785_/Y VGND VGND VPWR VPWR _12790_/Y sky130_fd_sc_hd__o21ai_1
X_11810_ _11810_/A _11810_/B VGND VGND VPWR VPWR _11810_/X sky130_fd_sc_hd__or2_1
XFILLER_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11771_/A _11741_/B VGND VGND VPWR VPWR _11741_/X sky130_fd_sc_hd__or2_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11672_ _14144_/A _11564_/B _11564_/Y _11566_/A VGND VGND VPWR VPWR _12643_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14457_/Y _14458_/Y _14459_/Y VGND VGND VPWR VPWR _14460_/X sky130_fd_sc_hd__o21a_1
XFILLER_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14391_ _15605_/A _14389_/X _14390_/X VGND VGND VPWR VPWR _14391_/X sky130_fd_sc_hd__o21a_1
X_13411_ _13411_/A VGND VGND VPWR VPWR _13411_/Y sky130_fd_sc_hd__inv_2
X_10623_ _10623_/A _12919_/A VGND VGND VPWR VPWR _12041_/A sky130_fd_sc_hd__or2_1
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16130_ _16243_/A VGND VGND VPWR VPWR _16205_/A sky130_fd_sc_hd__clkbuf_2
X_13342_ _14039_/A VGND VGND VPWR VPWR _15467_/A sky130_fd_sc_hd__buf_1
X_10554_ _11854_/A _10554_/B VGND VGND VPWR VPWR _10554_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16061_ _16123_/A _16123_/B VGND VGND VPWR VPWR _16061_/X sky130_fd_sc_hd__and2_1
X_13273_ _14722_/A _13272_/B _11413_/X _13272_/Y VGND VGND VPWR VPWR _13273_/X sky130_fd_sc_hd__o2bb2a_1
X_10485_ _12930_/A VGND VGND VPWR VPWR _11841_/A sky130_fd_sc_hd__inv_2
XFILLER_108_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12224_ _12224_/A _12224_/B VGND VGND VPWR VPWR _12224_/Y sky130_fd_sc_hd__nand2_1
X_15012_ _15042_/A _15042_/B VGND VGND VPWR VPWR _15061_/A sky130_fd_sc_hd__and2_1
XFILLER_6_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12155_ _13200_/A _12155_/B VGND VGND VPWR VPWR _12155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11106_ _11106_/A VGND VGND VPWR VPWR _11106_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12086_ _12087_/A _12087_/B VGND VGND VPWR VPWR _12088_/A sky130_fd_sc_hd__and2_1
X_15914_ _15909_/Y _15913_/Y _15909_/Y _15913_/Y VGND VGND VPWR VPWR _15972_/B sky130_fd_sc_hd__a2bb2o_1
X_11037_ _15075_/A VGND VGND VPWR VPWR _13918_/A sky130_fd_sc_hd__buf_1
XFILLER_77_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15845_ _14208_/A _15844_/X _12625_/X VGND VGND VPWR VPWR _15845_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15776_ _15774_/Y _15775_/X _15774_/Y _15775_/X VGND VGND VPWR VPWR _15782_/B sky130_fd_sc_hd__o2bb2a_1
X_12988_ _12929_/X _12987_/Y _12929_/X _12987_/Y VGND VGND VPWR VPWR _13018_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14727_ _14727_/A _14727_/B VGND VGND VPWR VPWR _14727_/X sky130_fd_sc_hd__or2_1
X_11939_ _11939_/A _11976_/B VGND VGND VPWR VPWR _11939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14658_ _15343_/A _14658_/B VGND VGND VPWR VPWR _14658_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13609_ _13609_/A _13609_/B VGND VGND VPWR VPWR _13609_/X sky130_fd_sc_hd__and2_1
XFILLER_20_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16328_ _16328_/A _16328_/B VGND VGND VPWR VPWR _16328_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14589_ _14539_/Y _14587_/X _14588_/Y VGND VGND VPWR VPWR _14589_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16259_ _16202_/Y _16256_/X _16258_/Y VGND VGND VPWR VPWR _16259_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09702_ _09695_/A _09695_/B _09698_/A VGND VGND VPWR VPWR _09970_/A sky130_fd_sc_hd__a21bo_1
XFILLER_95_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09633_ _08679_/A _09028_/A _09540_/X VGND VGND VPWR VPWR _09633_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_82_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09564_ _09478_/A _09518_/B _09478_/A _09518_/B VGND VGND VPWR VPWR _09564_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08515_ _09561_/A _08989_/A _08514_/Y VGND VGND VPWR VPWR _08515_/X sky130_fd_sc_hd__a21o_1
X_09495_ _08814_/X _09465_/X _08814_/X _09465_/X VGND VGND VPWR VPWR _09496_/B sky130_fd_sc_hd__o2bb2a_1
X_08446_ _08446_/A VGND VGND VPWR VPWR _08446_/Y sky130_fd_sc_hd__inv_2
X_08377_ _08242_/A input6/X _08307_/B _08460_/A VGND VGND VPWR VPWR _08465_/A sky130_fd_sc_hd__o22a_1
XFILLER_11_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10270_ _11742_/A VGND VGND VPWR VPWR _10325_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13960_ _15418_/A _13960_/B VGND VGND VPWR VPWR _13960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12911_ _12923_/A _12924_/B VGND VGND VPWR VPWR _12911_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15630_ _15673_/A _15673_/B VGND VGND VPWR VPWR _15630_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13891_ _14745_/A _13860_/B _13860_/Y VGND VGND VPWR VPWR _13891_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12842_ _12842_/A _12842_/B VGND VGND VPWR VPWR _12842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12773_/A _12773_/B VGND VGND VPWR VPWR _12773_/Y sky130_fd_sc_hd__nand2_1
X_15561_ _12425_/A _12426_/B _15560_/Y _15161_/A VGND VGND VPWR VPWR _15561_/X sky130_fd_sc_hd__o22a_1
XFILLER_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15492_ _15440_/A _15440_/B _15440_/A _15440_/B VGND VGND VPWR VPWR _15492_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _15208_/A _14512_/B VGND VGND VPWR VPWR _14512_/X sky130_fd_sc_hd__or2_1
X_11724_ _11724_/A _11730_/A VGND VGND VPWR VPWR _11724_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11655_/A _11654_/X VGND VGND VPWR VPWR _11655_/X sky130_fd_sc_hd__or2b_1
X_14443_ _14421_/A _14421_/B _14421_/Y VGND VGND VPWR VPWR _14443_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14374_ _14248_/A _14371_/X _14373_/Y _14249_/B _14373_/A VGND VGND VPWR VPWR _14375_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10606_ _10744_/A _10632_/B VGND VGND VPWR VPWR _10606_/Y sky130_fd_sc_hd__nor2_1
X_11586_ _09667_/Y _11585_/Y _09667_/Y _11585_/Y VGND VGND VPWR VPWR _11587_/B sky130_fd_sc_hd__o2bb2a_1
X_16113_ _16070_/X _16111_/X _16163_/B VGND VGND VPWR VPWR _16113_/X sky130_fd_sc_hd__o21a_1
X_13325_ _13365_/A _13365_/B VGND VGND VPWR VPWR _13388_/A sky130_fd_sc_hd__and2_1
X_10537_ _12934_/A VGND VGND VPWR VPWR _11867_/A sky130_fd_sc_hd__inv_2
XFILLER_6_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16044_ _16044_/A _16044_/B VGND VGND VPWR VPWR _16044_/Y sky130_fd_sc_hd__nand2_1
X_13256_ _15078_/A VGND VGND VPWR VPWR _14425_/A sky130_fd_sc_hd__inv_2
X_10468_ _10454_/X _10467_/Y _10454_/X _10467_/Y VGND VGND VPWR VPWR _10552_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ _12207_/A _12151_/X VGND VGND VPWR VPWR _12207_/X sky130_fd_sc_hd__or2b_1
XFILLER_97_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13187_ _13174_/Y _13185_/X _13186_/Y VGND VGND VPWR VPWR _13187_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10399_ _10359_/X _10398_/X _10359_/X _10398_/X VGND VGND VPWR VPWR _10400_/B sky130_fd_sc_hd__a2bb2o_1
X_12138_ _12228_/A _12136_/X _12137_/X VGND VGND VPWR VPWR _12138_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12069_ _12069_/A VGND VGND VPWR VPWR _12069_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15828_ _15826_/Y _15827_/X _15826_/Y _15827_/X VGND VGND VPWR VPWR _15828_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_80_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15759_ _16101_/A VGND VGND VPWR VPWR _16104_/A sky130_fd_sc_hd__buf_1
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09280_ _08623_/A _09802_/A _09224_/A VGND VGND VPWR VPWR _09280_/X sky130_fd_sc_hd__o21a_1
X_08300_ _08298_/X _08299_/X _08298_/A _08299_/X VGND VGND VPWR VPWR _08400_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08995_ _08990_/Y _08994_/X _08990_/Y _08994_/X VGND VGND VPWR VPWR _08995_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09616_ _09498_/A _09498_/B _09498_/Y VGND VGND VPWR VPWR _09616_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09547_ _09547_/A _09547_/B VGND VGND VPWR VPWR _09648_/B sky130_fd_sc_hd__and2_1
XFILLER_70_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09478_ _09478_/A _09478_/B VGND VGND VPWR VPWR _09478_/X sky130_fd_sc_hd__or2_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08429_ _08429_/A VGND VGND VPWR VPWR _08429_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11440_ _15529_/A _11440_/B VGND VGND VPWR VPWR _11440_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11371_ _08896_/X _11371_/B VGND VGND VPWR VPWR _11371_/X sky130_fd_sc_hd__and2b_1
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14090_ _14050_/X _14089_/X _14050_/X _14089_/X VGND VGND VPWR VPWR _14090_/Y sky130_fd_sc_hd__a2bb2oi_1
X_13110_ _13082_/Y _13108_/X _13109_/Y VGND VGND VPWR VPWR _13110_/X sky130_fd_sc_hd__o21a_1
X_10322_ _10344_/B _10322_/B VGND VGND VPWR VPWR _11776_/A sky130_fd_sc_hd__or2_1
XFILLER_125_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13041_ _15234_/A _13125_/B VGND VGND VPWR VPWR _13041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10253_ _10250_/Y _10251_/Y _10252_/Y VGND VGND VPWR VPWR _10254_/B sky130_fd_sc_hd__o21ai_2
XFILLER_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10184_ _10251_/A _10170_/B _10170_/Y _10377_/A VGND VGND VPWR VPWR _10462_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14992_ _14975_/X _14991_/X _14975_/X _14991_/X VGND VGND VPWR VPWR _15778_/B sky130_fd_sc_hd__a2bb2oi_4
XFILLER_59_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13943_ _13929_/Y _13941_/Y _13942_/Y VGND VGND VPWR VPWR _13943_/X sky130_fd_sc_hd__o21a_1
XFILLER_47_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13874_ _13874_/A _13874_/B VGND VGND VPWR VPWR _13874_/X sky130_fd_sc_hd__or2_1
XFILLER_47_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15613_ _14387_/X _15612_/X _14387_/X _15612_/X VGND VGND VPWR VPWR _15677_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12825_ _12825_/A _12838_/B VGND VGND VPWR VPWR _12825_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15544_ _15544_/A _15544_/B VGND VGND VPWR VPWR _15593_/B sky130_fd_sc_hd__or2_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12756_ _12765_/A _12765_/B VGND VGND VPWR VPWR _12756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11707_ _11707_/A VGND VGND VPWR VPWR _11707_/X sky130_fd_sc_hd__clkbuf_2
X_15475_ _15470_/A _15470_/B _15470_/Y _15474_/X VGND VGND VPWR VPWR _15475_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _10978_/A _12670_/A _10978_/Y _12670_/Y VGND VGND VPWR VPWR _12688_/B sky130_fd_sc_hd__o22a_1
X_11638_ _12387_/A _11638_/B VGND VGND VPWR VPWR _11638_/Y sky130_fd_sc_hd__nor2_1
X_14426_ _11778_/Y _14416_/A _11778_/Y _14416_/A VGND VGND VPWR VPWR _14427_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_128_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14357_ _14906_/A _13408_/B _13408_/X VGND VGND VPWR VPWR _14358_/A sky130_fd_sc_hd__o21ba_1
XFILLER_7_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11569_ _11569_/A _11569_/B VGND VGND VPWR VPWR _14149_/A sky130_fd_sc_hd__or2_1
X_13308_ _13210_/Y _13307_/X _13210_/Y _13307_/X VGND VGND VPWR VPWR _13309_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14288_ _15910_/A _14288_/B VGND VGND VPWR VPWR _14288_/X sky130_fd_sc_hd__or2_1
X_16027_ _16027_/A _16027_/B VGND VGND VPWR VPWR _16027_/Y sky130_fd_sc_hd__nand2_1
X_13239_ _13195_/X _13238_/Y _13195_/X _13238_/Y VGND VGND VPWR VPWR _13291_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08780_ _09333_/A _09472_/B _08711_/Y VGND VGND VPWR VPWR _08781_/A sky130_fd_sc_hd__a21oi_2
XFILLER_84_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09401_ _09401_/A _09707_/B VGND VGND VPWR VPWR _09401_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09332_ _09332_/A _10132_/A VGND VGND VPWR VPWR _10038_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09263_ _09263_/A _09263_/B VGND VGND VPWR VPWR _09263_/X sky130_fd_sc_hd__or2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09194_ _09341_/A _09161_/Y _09342_/A VGND VGND VPWR VPWR _09194_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08978_ _08978_/A _08978_/B VGND VGND VPWR VPWR _11364_/B sky130_fd_sc_hd__or2_1
XFILLER_29_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10940_ _10940_/A VGND VGND VPWR VPWR _11590_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12610_ _12610_/A VGND VGND VPWR VPWR _12610_/Y sky130_fd_sc_hd__inv_2
X_10871_ _12055_/A VGND VGND VPWR VPWR _10875_/A sky130_fd_sc_hd__inv_2
XFILLER_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13590_ _13637_/A _13638_/B VGND VGND VPWR VPWR _13590_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12541_ _12541_/A _12541_/B VGND VGND VPWR VPWR _12541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15260_ _15219_/X _15259_/Y _15219_/X _15259_/Y VGND VGND VPWR VPWR _15261_/B sky130_fd_sc_hd__a2bb2o_1
X_12472_ _12442_/Y _12471_/X _12442_/Y _12471_/X VGND VGND VPWR VPWR _12472_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14211_ _14101_/A _14101_/B _14101_/Y VGND VGND VPWR VPWR _14211_/X sky130_fd_sc_hd__o21a_1
X_11423_ _13349_/A _11242_/B _11242_/Y VGND VGND VPWR VPWR _11423_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15191_ _15125_/A _15125_/B _15125_/Y VGND VGND VPWR VPWR _15191_/Y sky130_fd_sc_hd__o21ai_1
X_11354_ _14064_/A _11353_/B _11353_/Y VGND VGND VPWR VPWR _11354_/Y sky130_fd_sc_hd__o21ai_1
X_14142_ _14065_/X _14141_/X _14065_/X _14141_/X VGND VGND VPWR VPWR _14145_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14073_ _14000_/Y _14072_/X _14000_/Y _14072_/X VGND VGND VPWR VPWR _14073_/X sky130_fd_sc_hd__a2bb2o_1
X_11285_ _09663_/X _11284_/X _09663_/X _11284_/X VGND VGND VPWR VPWR _11286_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_3_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10305_ _10305_/A VGND VGND VPWR VPWR _10305_/Y sky130_fd_sc_hd__inv_2
X_13024_ _14412_/A _13024_/B VGND VGND VPWR VPWR _13024_/X sky130_fd_sc_hd__or2_1
X_10236_ _10234_/Y _10235_/X _10175_/Y VGND VGND VPWR VPWR _10236_/Y sky130_fd_sc_hd__o21ai_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10167_ _10167_/A _10167_/B VGND VGND VPWR VPWR _10167_/Y sky130_fd_sc_hd__nor2_1
X_14975_ _14970_/Y _14974_/X _14970_/Y _14974_/X VGND VGND VPWR VPWR _14975_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_47_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10098_ _10098_/A _10098_/B VGND VGND VPWR VPWR _10099_/A sky130_fd_sc_hd__or2_1
X_13926_ _13926_/A VGND VGND VPWR VPWR _15400_/A sky130_fd_sc_hd__buf_1
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13857_ _13806_/Y _13855_/X _13856_/Y VGND VGND VPWR VPWR _13857_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13788_ _13783_/X _13787_/Y _13783_/X _13787_/Y VGND VGND VPWR VPWR _13865_/B sky130_fd_sc_hd__a2bb2o_1
X_12808_ _12773_/A _12773_/B _12773_/Y VGND VGND VPWR VPWR _12808_/Y sky130_fd_sc_hd__o21ai_1
X_15527_ _15461_/A _15461_/B _15461_/Y VGND VGND VPWR VPWR _15527_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12739_ _12692_/A _12692_/B _12692_/Y VGND VGND VPWR VPWR _12739_/X sky130_fd_sc_hd__a21o_1
X_15458_ _15458_/A _15458_/B VGND VGND VPWR VPWR _15458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14409_ _15440_/A VGND VGND VPWR VPWR _14774_/A sky130_fd_sc_hd__buf_1
XFILLER_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15389_ _15400_/A _15400_/B VGND VGND VPWR VPWR _15465_/A sky130_fd_sc_hd__and2_1
XFILLER_128_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09950_ _11770_/A VGND VGND VPWR VPWR _13560_/A sky130_fd_sc_hd__buf_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08901_ _08974_/A _08974_/B VGND VGND VPWR VPWR _08901_/X sky130_fd_sc_hd__and2_1
XFILLER_97_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09865_/X _08806_/Y _09865_/X _08806_/Y VGND VGND VPWR VPWR _09882_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _08831_/X _08725_/Y _08831_/A _08725_/Y VGND VGND VPWR VPWR _08834_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08763_ _09332_/A VGND VGND VPWR VPWR _09484_/A sky130_fd_sc_hd__buf_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08694_ _08694_/A _10120_/B VGND VGND VPWR VPWR _08871_/B sky130_fd_sc_hd__and2_1
XFILLER_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09315_ _09275_/A _09275_/B _09275_/X _10541_/A VGND VGND VPWR VPWR _10660_/A sky130_fd_sc_hd__a22o_1
X_09246_ _08572_/A _09858_/A _09318_/A VGND VGND VPWR VPWR _09246_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09177_ _09431_/A _09180_/B VGND VGND VPWR VPWR _09177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11070_ _12047_/A _10907_/B _10907_/Y VGND VGND VPWR VPWR _11070_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10021_ _09458_/A _10124_/A _10061_/B _10020_/X VGND VGND VPWR VPWR _10021_/X sky130_fd_sc_hd__o22a_1
XFILLER_130_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14760_ _15181_/A _14761_/B VGND VGND VPWR VPWR _14762_/A sky130_fd_sc_hd__and2_1
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11972_ _13073_/A _11972_/B VGND VGND VPWR VPWR _11972_/Y sky130_fd_sc_hd__nand2_1
X_13711_ _15046_/A _13504_/B _13504_/Y VGND VGND VPWR VPWR _13711_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10923_ _11011_/A _10920_/X _10922_/X VGND VGND VPWR VPWR _10923_/X sky130_fd_sc_hd__o21a_1
X_14691_ _15347_/A _14662_/B _14662_/Y VGND VGND VPWR VPWR _14691_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16430_ _16416_/Y _16447_/B _16428_/Y _16415_/X _16429_/X VGND VGND VPWR VPWR _16445_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_72_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13642_ _15122_/A _13642_/B VGND VGND VPWR VPWR _13642_/Y sky130_fd_sc_hd__nand2_1
X_10854_ _10854_/A VGND VGND VPWR VPWR _10854_/Y sky130_fd_sc_hd__inv_2
X_16361_ _16361_/A VGND VGND VPWR VPWR _16361_/X sky130_fd_sc_hd__buf_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _12135_/A _12914_/B _12916_/A _12914_/Y VGND VGND VPWR VPWR _13573_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12524_ _13442_/A _12306_/B _12306_/Y VGND VGND VPWR VPWR _12525_/B sky130_fd_sc_hd__o21a_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ _14582_/A _15255_/B _15255_/Y VGND VGND VPWR VPWR _15312_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10785_ _10785_/A VGND VGND VPWR VPWR _10785_/Y sky130_fd_sc_hd__inv_2
X_16292_ _16263_/X _16291_/Y _16263_/X _16291_/Y VGND VGND VPWR VPWR _16330_/B sky130_fd_sc_hd__o2bb2a_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15243_ _15243_/A _15243_/B VGND VGND VPWR VPWR _15243_/Y sky130_fd_sc_hd__nand2_1
X_12455_ _12454_/Y _12364_/X _12390_/Y VGND VGND VPWR VPWR _12480_/A sky130_fd_sc_hd__o21ai_2
XFILLER_125_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15174_ _15556_/A _15556_/B VGND VGND VPWR VPWR _15174_/Y sky130_fd_sc_hd__nand2_1
X_12386_ _12368_/X _12385_/X _12368_/X _12385_/X VGND VGND VPWR VPWR _12449_/B sky130_fd_sc_hd__a2bb2o_1
X_11406_ _08942_/A _08942_/B _08942_/Y VGND VGND VPWR VPWR _11407_/A sky130_fd_sc_hd__o21ai_1
XFILLER_126_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14125_ _14126_/A _14127_/A VGND VGND VPWR VPWR _14125_/Y sky130_fd_sc_hd__nor2_1
X_11337_ _11303_/X _11336_/X _11303_/X _11336_/X VGND VGND VPWR VPWR _11498_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14056_ _14056_/A _14056_/B VGND VGND VPWR VPWR _14056_/X sky130_fd_sc_hd__or2_1
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11268_ _09431_/B _09377_/B _09377_/X VGND VGND VPWR VPWR _11269_/B sky130_fd_sc_hd__a21boi_1
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13007_ _13007_/A VGND VGND VPWR VPWR _13007_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10219_ _10455_/A _11231_/A VGND VGND VPWR VPWR _11745_/A sky130_fd_sc_hd__or2_1
X_11199_ _11199_/A VGND VGND VPWR VPWR _11199_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14958_ _15353_/A _14958_/B VGND VGND VPWR VPWR _14958_/Y sky130_fd_sc_hd__nor2_1
X_14889_ _15534_/A _14914_/B VGND VGND VPWR VPWR _14889_/Y sky130_fd_sc_hd__nor2_1
X_13909_ _15410_/A _13952_/B VGND VGND VPWR VPWR _13909_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09100_ _09709_/A VGND VGND VPWR VPWR _09407_/A sky130_fd_sc_hd__buf_1
X_09031_ _09538_/B _09031_/B VGND VGND VPWR VPWR _09032_/B sky130_fd_sc_hd__or2_1
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09933_ _09932_/A _09932_/B _09932_/X VGND VGND VPWR VPWR _09933_/X sky130_fd_sc_hd__a21bo_1
X_09864_ _09863_/A _09863_/B _09863_/X VGND VGND VPWR VPWR _09864_/X sky130_fd_sc_hd__a21bo_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _08814_/X _08727_/X _08814_/A _08727_/X VGND VGND VPWR VPWR _08817_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09795_ _09196_/Y _09794_/A _09198_/X _09794_/Y VGND VGND VPWR VPWR _10618_/A sky130_fd_sc_hd__o22a_4
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08746_ _10008_/A _09448_/B VGND VGND VPWR VPWR _08746_/X sky130_fd_sc_hd__or2_1
XFILLER_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08677_ _09235_/A _08677_/B VGND VGND VPWR VPWR _08678_/A sky130_fd_sc_hd__or2_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10570_ _10569_/A _10569_/B _10569_/Y _10982_/A VGND VGND VPWR VPWR _11918_/A sky130_fd_sc_hd__o211a_1
X_09229_ _09800_/A VGND VGND VPWR VPWR _09687_/A sky130_fd_sc_hd__inv_2
XFILLER_107_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12240_ _14036_/A _12224_/B _12224_/Y _12239_/X VGND VGND VPWR VPWR _12240_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12171_ _12261_/A VGND VGND VPWR VPWR _12781_/A sky130_fd_sc_hd__buf_1
XFILLER_107_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11122_ _12095_/A _11122_/B VGND VGND VPWR VPWR _11122_/Y sky130_fd_sc_hd__nor2_1
X_15930_ _15958_/A _15958_/B VGND VGND VPWR VPWR _16008_/A sky130_fd_sc_hd__and2_1
XFILLER_89_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11053_ _12825_/A VGND VGND VPWR VPWR _15084_/A sky130_fd_sc_hd__buf_1
XFILLER_49_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15861_ _14190_/X _15847_/X _14190_/X _15847_/X VGND VGND VPWR VPWR _15900_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10004_ _10344_/B VGND VGND VPWR VPWR _10446_/A sky130_fd_sc_hd__inv_2
X_14812_ _14812_/A _14812_/B VGND VGND VPWR VPWR _14812_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15792_ _15668_/Y _15791_/Y _15668_/Y _15791_/Y VGND VGND VPWR VPWR _16227_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14743_ _15349_/A _14743_/B VGND VGND VPWR VPWR _14743_/Y sky130_fd_sc_hd__nor2_1
X_11955_ _11892_/A _11892_/B _11892_/Y VGND VGND VPWR VPWR _11955_/Y sky130_fd_sc_hd__o21ai_1
X_10906_ _10906_/A VGND VGND VPWR VPWR _11065_/A sky130_fd_sc_hd__inv_2
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14674_ _14674_/A _14674_/B VGND VGND VPWR VPWR _14674_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16413_ _16474_/Q VGND VGND VPWR VPWR _16437_/D sky130_fd_sc_hd__inv_2
X_11886_ _11886_/A _12041_/A VGND VGND VPWR VPWR _11959_/A sky130_fd_sc_hd__or2_1
X_13625_ _13625_/A VGND VGND VPWR VPWR _15134_/A sky130_fd_sc_hd__buf_1
XFILLER_32_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10837_ _12005_/A _10944_/B _10836_/Y VGND VGND VPWR VPWR _10837_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16344_ _08230_/X _16470_/Q _08233_/X _16392_/A _16343_/X VGND VGND VPWR VPWR _16470_/D
+ sky130_fd_sc_hd__o221a_2
X_10768_ _11964_/A VGND VGND VPWR VPWR _14564_/A sky130_fd_sc_hd__buf_1
XFILLER_80_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13556_ _13556_/A _13556_/B VGND VGND VPWR VPWR _13557_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16275_ _16137_/Y _16274_/Y _16137_/Y _16274_/Y VGND VGND VPWR VPWR _16277_/B sky130_fd_sc_hd__a2bb2o_1
X_12507_ _12506_/A _12506_/B _12506_/Y _11707_/X VGND VGND VPWR VPWR _12637_/A sky130_fd_sc_hd__o211a_1
X_13487_ _10669_/Y _11859_/A _10572_/Y _13486_/X VGND VGND VPWR VPWR _13487_/X sky130_fd_sc_hd__o22a_1
X_15226_ _15187_/A _15187_/B _15187_/Y _15225_/X VGND VGND VPWR VPWR _15226_/X sky130_fd_sc_hd__a2bb2o_1
X_10699_ _11933_/A _10789_/B _10698_/Y VGND VGND VPWR VPWR _10699_/Y sky130_fd_sc_hd__o21ai_1
X_12438_ _12437_/A _12437_/B _12437_/X VGND VGND VPWR VPWR _12439_/B sky130_fd_sc_hd__a21bo_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15157_ _15116_/A _15116_/B _15116_/Y _15156_/X VGND VGND VPWR VPWR _15157_/X sky130_fd_sc_hd__a2bb2o_1
X_12369_ _12369_/A _12369_/B VGND VGND VPWR VPWR _12369_/X sky130_fd_sc_hd__or2_1
XFILLER_114_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14108_ _14108_/A _14112_/B VGND VGND VPWR VPWR _14108_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15088_ _12835_/X _15144_/A _15087_/X VGND VGND VPWR VPWR _15088_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14039_ _14039_/A _14039_/B VGND VGND VPWR VPWR _14039_/X sky130_fd_sc_hd__and2_1
XFILLER_67_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08600_ _08599_/A _08348_/Y _08599_/Y _08348_/A VGND VGND VPWR VPWR _08601_/B sky130_fd_sc_hd__o22a_1
XFILLER_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09580_ _09486_/A _09486_/B _09486_/Y VGND VGND VPWR VPWR _09580_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08531_ _09474_/B VGND VGND VPWR VPWR _08692_/A sky130_fd_sc_hd__buf_1
X_08462_ _08697_/A VGND VGND VPWR VPWR _09448_/A sky130_fd_sc_hd__inv_2
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08393_ _08393_/A1 input18/X _08392_/A _08399_/A _08392_/Y VGND VGND VPWR VPWR _08394_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09014_ _09488_/A _09020_/S _08565_/B VGND VGND VPWR VPWR _09014_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09916_ _10947_/A _10946_/A VGND VGND VPWR VPWR _09916_/X sky130_fd_sc_hd__or2_1
XFILLER_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09847_ _10491_/A _09846_/X VGND VGND VPWR VPWR _09848_/B sky130_fd_sc_hd__or2b_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09778_ _09779_/A _09779_/B VGND VGND VPWR VPWR _09778_/Y sky130_fd_sc_hd__nor2_1
X_08729_ _08729_/A VGND VGND VPWR VPWR _08729_/Y sky130_fd_sc_hd__inv_2
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11776_/A _11728_/B _11728_/X _11739_/Y VGND VGND VPWR VPWR _11741_/B sky130_fd_sc_hd__a22o_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11671_ _15554_/A _11673_/B VGND VGND VPWR VPWR _11671_/X sky130_fd_sc_hd__and2_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14390_ _15960_/A _14390_/B VGND VGND VPWR VPWR _14390_/X sky130_fd_sc_hd__or2_1
X_13410_ _13356_/Y _13409_/X _13356_/Y _13409_/X VGND VGND VPWR VPWR _13411_/A sky130_fd_sc_hd__a2bb2o_1
X_10622_ _10622_/A _12916_/A _10622_/C VGND VGND VPWR VPWR _12919_/A sky130_fd_sc_hd__and3_1
XFILLER_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13341_ _13341_/A VGND VGND VPWR VPWR _14039_/A sky130_fd_sc_hd__buf_1
X_10553_ _10550_/Y _12696_/A _10452_/X _10552_/Y VGND VGND VPWR VPWR _10553_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16060_ _16054_/X _16059_/X _16054_/X _16059_/X VGND VGND VPWR VPWR _16123_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13272_ _15087_/A _13272_/B VGND VGND VPWR VPWR _13272_/Y sky130_fd_sc_hd__nor2_1
X_15011_ _11998_/X _15004_/X _11998_/X _15004_/X VGND VGND VPWR VPWR _15042_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10484_ _09849_/Y _10483_/X _09851_/A _09850_/Y _10792_/A VGND VGND VPWR VPWR _12930_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12223_ _12140_/X _12222_/X _12140_/X _12222_/X VGND VGND VPWR VPWR _12224_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12154_ _12204_/A _12152_/X _12153_/X VGND VGND VPWR VPWR _12154_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11105_ _11105_/A VGND VGND VPWR VPWR _11105_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12085_ _10978_/A _12084_/A _10978_/Y _12174_/B VGND VGND VPWR VPWR _12087_/B sky130_fd_sc_hd__o22a_1
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15913_ _15978_/A _15978_/B _15912_/Y VGND VGND VPWR VPWR _15913_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11036_ _12844_/A VGND VGND VPWR VPWR _15075_/A sky130_fd_sc_hd__clkbuf_2
X_15844_ _14214_/A _15843_/X _12623_/X VGND VGND VPWR VPWR _15844_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15775_ _15665_/X _15775_/B VGND VGND VPWR VPWR _15775_/X sky130_fd_sc_hd__and2b_1
XFILLER_92_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14726_ _14807_/A _14724_/X _14807_/B VGND VGND VPWR VPWR _14726_/Y sky130_fd_sc_hd__o21bai_1
X_12987_ _14465_/A _12930_/B _12930_/Y VGND VGND VPWR VPWR _12987_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11938_ _11979_/A _11937_/Y _11979_/A _11937_/Y VGND VGND VPWR VPWR _11976_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14657_ _14622_/Y _14655_/X _14656_/Y VGND VGND VPWR VPWR _14657_/X sky130_fd_sc_hd__o21a_1
X_11869_ _11844_/X _11868_/Y _11844_/X _11868_/Y VGND VGND VPWR VPWR _11907_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14588_ _14588_/A _14588_/B VGND VGND VPWR VPWR _14588_/Y sky130_fd_sc_hd__nand2_1
X_13608_ _13573_/X _13607_/X _13573_/X _13607_/X VGND VGND VPWR VPWR _13609_/B sky130_fd_sc_hd__a2bb2o_1
X_16327_ _16299_/Y _16325_/X _16326_/Y VGND VGND VPWR VPWR _16327_/X sky130_fd_sc_hd__o21a_1
X_13539_ _15042_/A _13510_/B _13510_/Y _13538_/X VGND VGND VPWR VPWR _13539_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16258_ _16324_/A _16258_/B VGND VGND VPWR VPWR _16258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16189_ _16189_/A _16189_/B VGND VGND VPWR VPWR _16260_/A sky130_fd_sc_hd__or2_1
XFILLER_114_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15209_ _15143_/A _15143_/B _15143_/Y VGND VGND VPWR VPWR _15209_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09701_ _09701_/A VGND VGND VPWR VPWR _09770_/A sky130_fd_sc_hd__inv_2
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09632_ _09632_/A VGND VGND VPWR VPWR _09632_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09563_ _09563_/A VGND VGND VPWR VPWR _09563_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08514_ _09561_/A _08989_/A VGND VGND VPWR VPWR _08514_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09494_ _09494_/A _09494_/B VGND VGND VPWR VPWR _09494_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08445_ _08555_/B _08439_/Y _09333_/A VGND VGND VPWR VPWR _08446_/A sky130_fd_sc_hd__o21ai_1
XFILLER_24_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08376_ input5/X _08245_/B _08312_/B _08454_/A VGND VGND VPWR VPWR _08460_/A sky130_fd_sc_hd__o22a_1
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13890_ _13890_/A VGND VGND VPWR VPWR _15418_/A sky130_fd_sc_hd__buf_1
XFILLER_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12910_ _12837_/X _12909_/Y _12837_/X _12909_/Y VGND VGND VPWR VPWR _12924_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_104_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12841_ _12822_/Y _12839_/X _12840_/Y VGND VGND VPWR VPWR _12841_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12772_ _12747_/Y _12770_/X _12771_/Y VGND VGND VPWR VPWR _12772_/X sky130_fd_sc_hd__o21a_1
X_15560_ _15560_/A VGND VGND VPWR VPWR _15560_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15491_ _15552_/A _15552_/B VGND VGND VPWR VPWR _15491_/X sky130_fd_sc_hd__and2_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14565_/A _14509_/X _14510_/X VGND VGND VPWR VPWR _14511_/X sky130_fd_sc_hd__o21a_1
X_11723_ _12704_/A _11733_/B _12704_/A _11733_/B VGND VGND VPWR VPWR _11730_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _13989_/A _11654_/B VGND VGND VPWR VPWR _11654_/X sky130_fd_sc_hd__or2_1
X_14442_ _14469_/A _14469_/B VGND VGND VPWR VPWR _14442_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10605_ _10526_/X _10604_/Y _10526_/X _10604_/Y VGND VGND VPWR VPWR _10632_/B sky130_fd_sc_hd__a2bb2o_1
X_14373_ _14373_/A VGND VGND VPWR VPWR _14373_/Y sky130_fd_sc_hd__inv_2
X_16112_ _16112_/A _16112_/B VGND VGND VPWR VPWR _16163_/B sky130_fd_sc_hd__or2_1
X_11585_ _09569_/A _09569_/B _09569_/Y VGND VGND VPWR VPWR _11585_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_128_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13324_ _13293_/A _13323_/Y _13293_/A _13323_/Y VGND VGND VPWR VPWR _13365_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10536_ _09899_/Y _10535_/X _09901_/A _09900_/Y _10792_/A VGND VGND VPWR VPWR _12934_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16043_ _16007_/Y _16041_/X _16042_/Y VGND VGND VPWR VPWR _16043_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13255_ _14729_/A _13282_/B VGND VGND VPWR VPWR _13255_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10467_ _10467_/A VGND VGND VPWR VPWR _10467_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12206_ _14015_/A _12206_/B VGND VGND VPWR VPWR _12206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13186_ _13825_/A _13186_/B VGND VGND VPWR VPWR _13186_/Y sky130_fd_sc_hd__nand2_1
X_10398_ _13525_/A _10319_/B _11710_/A _10319_/B VGND VGND VPWR VPWR _10398_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12137_ _12137_/A _12137_/B VGND VGND VPWR VPWR _12137_/X sky130_fd_sc_hd__or2_1
XFILLER_96_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12068_ _12068_/A _12068_/B VGND VGND VPWR VPWR _12068_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11019_ _10917_/X _11018_/X _10917_/X _11018_/X VGND VGND VPWR VPWR _11089_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15827_ _14167_/A _14289_/X _14166_/X VGND VGND VPWR VPWR _15827_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15758_ _15765_/A _15758_/B VGND VGND VPWR VPWR _16101_/A sky130_fd_sc_hd__or2_1
XFILLER_80_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15689_ _15694_/A _15694_/B VGND VGND VPWR VPWR _15689_/Y sky130_fd_sc_hd__nor2_1
X_14709_ _15335_/A _14650_/B _14650_/Y VGND VGND VPWR VPWR _14709_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08230_ _08230_/A VGND VGND VPWR VPWR _08230_/X sky130_fd_sc_hd__buf_1
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08994_ _08992_/X _08993_/Y _08992_/X _08993_/Y VGND VGND VPWR VPWR _08994_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09615_ _09978_/A _09652_/B VGND VGND VPWR VPWR _09615_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09546_ _09546_/A VGND VGND VPWR VPWR _09546_/Y sky130_fd_sc_hd__inv_2
X_09477_ _09449_/Y _09475_/X _09476_/X VGND VGND VPWR VPWR _09477_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08428_ _09213_/B _08423_/X _08794_/A VGND VGND VPWR VPWR _08428_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08359_ input9/X _08278_/A _08399_/A VGND VGND VPWR VPWR _08359_/X sky130_fd_sc_hd__a21o_1
X_11370_ _12306_/A _11370_/B VGND VGND VPWR VPWR _11370_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10321_ _10216_/X _10320_/Y _10216_/X _10320_/Y VGND VGND VPWR VPWR _10322_/B sky130_fd_sc_hd__o2bb2a_1
X_13040_ _13033_/X _13039_/X _13033_/X _13039_/X VGND VGND VPWR VPWR _13125_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10252_ _10252_/A _10252_/B VGND VGND VPWR VPWR _10252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10183_ _10248_/A _10173_/B _10173_/Y _10182_/Y VGND VGND VPWR VPWR _10377_/A sky130_fd_sc_hd__o2bb2a_1
X_14991_ _14988_/X _14990_/Y _14988_/X _14990_/Y VGND VGND VPWR VPWR _14991_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_115_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13942_ _15400_/A _13942_/B VGND VGND VPWR VPWR _13942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13873_ _13873_/A _13873_/B VGND VGND VPWR VPWR _13874_/B sky130_fd_sc_hd__nor2_1
X_15612_ _15612_/A _14388_/X VGND VGND VPWR VPWR _15612_/X sky130_fd_sc_hd__or2b_1
X_12824_ _12762_/Y _12823_/Y _12762_/Y _12823_/Y VGND VGND VPWR VPWR _12838_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15543_ _15600_/A _15602_/A _15542_/X VGND VGND VPWR VPWR _15543_/X sky130_fd_sc_hd__o21a_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12755_ _12709_/X _12754_/X _12709_/X _12754_/X VGND VGND VPWR VPWR _12765_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11706_ _11706_/A VGND VGND VPWR VPWR _11707_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _15473_/A _15473_/B _12235_/X _15473_/Y VGND VGND VPWR VPWR _15474_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12686_/A _12686_/B VGND VGND VPWR VPWR _12686_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14425_ _14425_/A _14425_/B VGND VGND VPWR VPWR _14425_/Y sky130_fd_sc_hd__nor2_1
X_11637_ _11637_/A _11636_/X VGND VGND VPWR VPWR _11637_/X sky130_fd_sc_hd__or2b_1
XFILLER_30_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14356_ _14250_/Y _14355_/Y _14250_/Y _14355_/Y VGND VGND VPWR VPWR _14378_/A sky130_fd_sc_hd__a2bb2o_1
X_11568_ _08985_/X _11567_/X _08985_/X _11567_/X VGND VGND VPWR VPWR _11569_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13307_ _13215_/Y _13305_/Y _13306_/Y VGND VGND VPWR VPWR _13307_/X sky130_fd_sc_hd__o21a_1
X_10519_ _10428_/X _10518_/X _10622_/A _10518_/X VGND VGND VPWR VPWR _10523_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16026_ _14371_/X _15665_/B _14371_/X _15665_/B VGND VGND VPWR VPWR _16027_/B sky130_fd_sc_hd__a2bb2o_1
X_14287_ _14399_/A _14285_/X _14286_/X VGND VGND VPWR VPWR _14287_/X sky130_fd_sc_hd__o21a_1
X_11499_ _11498_/Y _11296_/X _11338_/Y VGND VGND VPWR VPWR _11499_/X sky130_fd_sc_hd__o21a_1
X_13238_ _13196_/A _13196_/B _13196_/Y VGND VGND VPWR VPWR _13238_/Y sky130_fd_sc_hd__o21ai_1
X_13169_ _15261_/A _13107_/B _13107_/Y VGND VGND VPWR VPWR _13169_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09400_ _09717_/A VGND VGND VPWR VPWR _09412_/A sky130_fd_sc_hd__inv_2
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09331_ _09331_/A _09331_/B VGND VGND VPWR VPWR _10035_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09262_ _10242_/A VGND VGND VPWR VPWR _09263_/B sky130_fd_sc_hd__buf_1
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09193_ _09193_/A VGND VGND VPWR VPWR _09193_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08977_ _08896_/X _08975_/X _11371_/B VGND VGND VPWR VPWR _08977_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10870_ _09946_/A _10869_/A _09946_/Y _10869_/Y _09445_/A VGND VGND VPWR VPWR _12055_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_71_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09529_ _09529_/A _09529_/B VGND VGND VPWR VPWR _09530_/A sky130_fd_sc_hd__or2_1
XFILLER_101_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12540_ _13438_/A _12312_/B _12312_/Y VGND VGND VPWR VPWR _12541_/B sky130_fd_sc_hd__o21a_1
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12471_ _12469_/Y _12470_/Y _12469_/Y _12470_/Y VGND VGND VPWR VPWR _12471_/X sky130_fd_sc_hd__o2bb2a_1
X_14210_ _15869_/A _14263_/B VGND VGND VPWR VPWR _14210_/Y sky130_fd_sc_hd__nor2_1
X_11422_ _14084_/A _11422_/B VGND VGND VPWR VPWR _11422_/Y sky130_fd_sc_hd__nor2_1
X_15190_ _15190_/A _15190_/B VGND VGND VPWR VPWR _15190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14141_ _14141_/A _14066_/X VGND VGND VPWR VPWR _14141_/X sky130_fd_sc_hd__or2b_1
XFILLER_125_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11353_ _14064_/A _11353_/B VGND VGND VPWR VPWR _11353_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14072_ _14070_/X _14071_/X _14070_/X _14071_/X VGND VGND VPWR VPWR _14072_/X sky130_fd_sc_hd__a2bb2o_1
X_11284_ _09995_/A _09664_/B _09664_/Y VGND VGND VPWR VPWR _11284_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10304_ _10248_/A _10173_/B _10173_/Y VGND VGND VPWR VPWR _10305_/A sky130_fd_sc_hd__a21oi_1
XFILLER_112_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13023_ _13070_/A _13021_/X _13022_/X VGND VGND VPWR VPWR _13023_/X sky130_fd_sc_hd__o21a_1
X_10235_ _10235_/A _10235_/B VGND VGND VPWR VPWR _10235_/X sky130_fd_sc_hd__and2_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10166_ _10126_/A _10126_/B _10127_/B VGND VGND VPWR VPWR _10167_/B sky130_fd_sc_hd__a21bo_1
XFILLER_120_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14974_ _14972_/X _14973_/Y _14972_/X _14973_/Y VGND VGND VPWR VPWR _14974_/X sky130_fd_sc_hd__o2bb2a_1
X_10097_ _11733_/A VGND VGND VPWR VPWR _10213_/A sky130_fd_sc_hd__inv_2
X_13925_ _15402_/A _13944_/B VGND VGND VPWR VPWR _13925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13856_ _14410_/A _13856_/B VGND VGND VPWR VPWR _13856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12807_ _12850_/A _12850_/B VGND VGND VPWR VPWR _12807_/Y sky130_fd_sc_hd__nor2_1
X_10999_ _13053_/A _10998_/B _10998_/Y VGND VGND VPWR VPWR _10999_/Y sky130_fd_sc_hd__o21ai_1
X_13787_ _12858_/A _13786_/B _13868_/A VGND VGND VPWR VPWR _13787_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15526_ _15529_/A _15529_/B VGND VGND VPWR VPWR _15526_/Y sky130_fd_sc_hd__nor2_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12777_/A _12777_/B VGND VGND VPWR VPWR _12738_/Y sky130_fd_sc_hd__nor2_1
X_15457_ _15405_/X _15456_/X _15405_/X _15456_/X VGND VGND VPWR VPWR _15458_/B sky130_fd_sc_hd__a2bb2o_1
X_12669_ _10964_/Y _12668_/Y _10821_/Y VGND VGND VPWR VPWR _12670_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14408_ _14408_/A VGND VGND VPWR VPWR _15552_/A sky130_fd_sc_hd__buf_1
X_15388_ _15332_/X _15387_/X _15332_/X _15387_/X VGND VGND VPWR VPWR _15400_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14339_ _14101_/A _13426_/B _13426_/Y VGND VGND VPWR VPWR _14339_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16009_ _15957_/X _16008_/X _15957_/X _16008_/X VGND VGND VPWR VPWR _16040_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09866_/X _08797_/A _09866_/X _08797_/A VGND VGND VPWR VPWR _09883_/A sky130_fd_sc_hd__a2bb2o_1
X_08900_ _08899_/Y _08862_/X _08899_/Y _08862_/X VGND VGND VPWR VPWR _08974_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A VGND VGND VPWR VPWR _08831_/X sky130_fd_sc_hd__buf_1
XFILLER_58_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08762_/A _10133_/A VGND VGND VPWR VPWR _08762_/Y sky130_fd_sc_hd__nor2_1
X_08693_ _08876_/A _08691_/X _08876_/B VGND VGND VPWR VPWR _08693_/X sky130_fd_sc_hd__o21ba_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09314_ _10438_/A _09312_/Y _09313_/Y VGND VGND VPWR VPWR _10541_/A sky130_fd_sc_hd__o21ai_2
X_09245_ _09555_/A _09734_/A VGND VGND VPWR VPWR _09318_/A sky130_fd_sc_hd__or2_1
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09176_ _09175_/Y _09040_/Y _09143_/Y VGND VGND VPWR VPWR _09180_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10020_ _08844_/A _09070_/A _08944_/X _10019_/X VGND VGND VPWR VPWR _10020_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11971_ _11948_/Y _11969_/X _11970_/Y VGND VGND VPWR VPWR _11971_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10922_ _14611_/A _10922_/B VGND VGND VPWR VPWR _10922_/X sky130_fd_sc_hd__or2_1
XFILLER_72_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13710_ _12854_/A _13649_/B _13709_/Y _13646_/X VGND VGND VPWR VPWR _13710_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14690_ _14741_/A _14741_/B VGND VGND VPWR VPWR _14776_/A sky130_fd_sc_hd__and2_1
XFILLER_72_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13641_ _13641_/A VGND VGND VPWR VPWR _15122_/A sky130_fd_sc_hd__buf_1
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10853_ _09421_/A _09421_/B _09421_/Y VGND VGND VPWR VPWR _10854_/A sky130_fd_sc_hd__o21ai_1
X_16360_ _16329_/X _16359_/Y _16329_/X _16359_/Y VGND VGND VPWR VPWR _16407_/D sky130_fd_sc_hd__a2bb2o_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _14429_/A _13574_/B VGND VGND VPWR VPWR _13607_/A sky130_fd_sc_hd__and2_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10784_ _09776_/A _09776_/B _09776_/Y VGND VGND VPWR VPWR _10785_/A sky130_fd_sc_hd__o21ai_1
X_16291_ _16264_/A _16330_/A _16264_/Y VGND VGND VPWR VPWR _16291_/Y sky130_fd_sc_hd__o21ai_1
X_12523_ _12522_/A _12522_/B _12522_/Y _11707_/X VGND VGND VPWR VPWR _12633_/A sky130_fd_sc_hd__o211a_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15311_ _15341_/A _15341_/B VGND VGND VPWR VPWR _15375_/A sky130_fd_sc_hd__and2_1
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15242_ _15225_/X _15241_/Y _15225_/X _15241_/Y VGND VGND VPWR VPWR _15243_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12454_ _12953_/A _12454_/B VGND VGND VPWR VPWR _12454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15173_ _15159_/Y _15172_/Y _15159_/Y _15172_/Y VGND VGND VPWR VPWR _15556_/B sky130_fd_sc_hd__a2bb2o_1
X_12385_ _13872_/A _12440_/B _13872_/A _12440_/B VGND VGND VPWR VPWR _12385_/X sky130_fd_sc_hd__a2bb2o_1
X_11405_ _11405_/A VGND VGND VPWR VPWR _11405_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14124_ _14059_/X _14123_/X _14059_/X _14123_/X VGND VGND VPWR VPWR _14127_/A sky130_fd_sc_hd__a2bb2o_1
X_11336_ _13786_/A _11504_/B _13786_/A _11504_/B VGND VGND VPWR VPWR _11336_/X sky130_fd_sc_hd__a2bb2o_1
X_14055_ _14109_/A _14024_/B _14024_/X _14054_/X VGND VGND VPWR VPWR _14055_/X sky130_fd_sc_hd__o22a_1
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11267_ _11177_/A _11094_/X _11176_/X VGND VGND VPWR VPWR _11267_/X sky130_fd_sc_hd__o21a_1
X_13006_ _13006_/A VGND VGND VPWR VPWR _13007_/A sky130_fd_sc_hd__buf_1
XFILLER_79_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11198_ _09424_/A _09131_/B _09131_/Y VGND VGND VPWR VPWR _11199_/A sky130_fd_sc_hd__o21ai_1
X_10218_ _10216_/X _10217_/Y _10216_/X _10217_/Y VGND VGND VPWR VPWR _11231_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_121_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10149_ _10151_/A VGND VGND VPWR VPWR _10241_/B sky130_fd_sc_hd__buf_1
X_14957_ _14956_/A _14956_/B _14956_/Y VGND VGND VPWR VPWR _14957_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14888_ _14820_/X _14887_/X _14820_/X _14887_/X VGND VGND VPWR VPWR _14914_/B sky130_fd_sc_hd__a2bb2o_1
X_13908_ _13851_/X _13907_/Y _13851_/X _13907_/Y VGND VGND VPWR VPWR _13952_/B sky130_fd_sc_hd__a2bb2o_1
X_13839_ _10906_/A _13837_/Y _13838_/Y VGND VGND VPWR VPWR _13839_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15509_ _15509_/A _15509_/B VGND VGND VPWR VPWR _15510_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09030_ _09539_/B _09030_/B VGND VGND VPWR VPWR _09031_/B sky130_fd_sc_hd__or2_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09932_ _09932_/A _09932_/B VGND VGND VPWR VPWR _09932_/X sky130_fd_sc_hd__or2_1
XFILLER_131_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09863_ _09863_/A _09863_/B VGND VGND VPWR VPWR _09863_/X sky130_fd_sc_hd__or2_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08814_ _08814_/A VGND VGND VPWR VPWR _08814_/X sky130_fd_sc_hd__buf_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09794_/A VGND VGND VPWR VPWR _09794_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08745_ _08745_/A VGND VGND VPWR VPWR _08745_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08676_ _10098_/B VGND VGND VPWR VPWR _08677_/B sky130_fd_sc_hd__inv_2
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09228_ _09228_/A _09228_/B VGND VGND VPWR VPWR _09800_/A sky130_fd_sc_hd__or2_1
XFILLER_108_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09159_ _08709_/Y _09158_/Y _08743_/X VGND VGND VPWR VPWR _09160_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12170_ _12170_/A VGND VGND VPWR VPWR _12261_/A sky130_fd_sc_hd__inv_2
XFILLER_107_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11121_ _12254_/A VGND VGND VPWR VPWR _13720_/A sky130_fd_sc_hd__buf_1
XFILLER_1_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11052_ _14427_/A _11079_/B VGND VGND VPWR VPWR _11234_/A sky130_fd_sc_hd__and2_1
XFILLER_89_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15860_ _15860_/A VGND VGND VPWR VPWR _15900_/A sky130_fd_sc_hd__inv_2
XFILLER_103_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10003_ _10001_/X _10002_/X _10001_/X _10002_/X VGND VGND VPWR VPWR _10344_/B sky130_fd_sc_hd__o2bb2a_2
X_14811_ _14723_/X _14810_/X _14723_/X _14810_/X VGND VGND VPWR VPWR _14812_/B sky130_fd_sc_hd__a2bb2o_1
X_15791_ _15669_/A _15669_/B _15669_/Y VGND VGND VPWR VPWR _15791_/Y sky130_fd_sc_hd__o21ai_1
X_14742_ _14776_/A _14740_/X _14741_/X VGND VGND VPWR VPWR _14742_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11954_ _13088_/A _11966_/B VGND VGND VPWR VPWR _11954_/Y sky130_fd_sc_hd__nor2_1
X_10905_ _15212_/B _12041_/B VGND VGND VPWR VPWR _10906_/A sky130_fd_sc_hd__or2_1
X_11885_ _11892_/A _11892_/B VGND VGND VPWR VPWR _11885_/Y sky130_fd_sc_hd__nor2_1
X_14673_ _12183_/Y _14672_/X _12183_/Y _14672_/X VGND VGND VPWR VPWR _14674_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16412_ _16469_/Q VGND VGND VPWR VPWR _16412_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13624_ _13624_/A VGND VGND VPWR VPWR _13624_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10836_ _12005_/A _10944_/B VGND VGND VPWR VPWR _10836_/Y sky130_fd_sc_hd__nand2_1
X_16343_ _16343_/A VGND VGND VPWR VPWR _16343_/X sky130_fd_sc_hd__buf_1
X_10767_ _10901_/A _10765_/X _10766_/X VGND VGND VPWR VPWR _10767_/X sky130_fd_sc_hd__o21a_1
X_13555_ _13535_/X _13554_/Y _13535_/X _13554_/Y VGND VGND VPWR VPWR _13556_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16274_ _16145_/Y _16271_/X _16273_/Y VGND VGND VPWR VPWR _16274_/Y sky130_fd_sc_hd__o21ai_1
X_12506_ _12506_/A _12506_/B VGND VGND VPWR VPWR _12506_/Y sky130_fd_sc_hd__nand2_1
X_10698_ _11933_/A _10789_/B VGND VGND VPWR VPWR _10698_/Y sky130_fd_sc_hd__nand2_1
X_13486_ _10550_/Y _11810_/A _10475_/Y _13485_/X VGND VGND VPWR VPWR _13486_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15225_ _15190_/A _15190_/B _15190_/Y _15224_/X VGND VGND VPWR VPWR _15225_/X sky130_fd_sc_hd__a2bb2o_1
X_12437_ _12437_/A _12437_/B VGND VGND VPWR VPWR _12437_/X sky130_fd_sc_hd__or2_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15156_ _15119_/A _15119_/B _15119_/Y _15155_/X VGND VGND VPWR VPWR _15156_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14107_ _14103_/Y _14105_/Y _14106_/Y VGND VGND VPWR VPWR _14112_/B sky130_fd_sc_hd__o21ai_1
X_12368_ _11273_/A _12367_/B _12367_/X _12260_/X VGND VGND VPWR VPWR _12368_/X sky130_fd_sc_hd__o22a_1
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12299_ _12247_/X _12298_/Y _12247_/X _12298_/Y VGND VGND VPWR VPWR _12300_/B sky130_fd_sc_hd__a2bb2o_1
X_15087_ _15087_/A _15087_/B VGND VGND VPWR VPWR _15087_/X sky130_fd_sc_hd__or2_1
X_11319_ _11319_/A VGND VGND VPWR VPWR _11518_/A sky130_fd_sc_hd__inv_2
XFILLER_4_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14038_ _13941_/Y _14037_/X _13941_/Y _14037_/X VGND VGND VPWR VPWR _14039_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15989_ _15973_/X _15988_/X _15973_/X _15988_/X VGND VGND VPWR VPWR _15991_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08530_ _09527_/A VGND VGND VPWR VPWR _09474_/B sky130_fd_sc_hd__inv_2
X_08461_ _08460_/A _08308_/Y _08460_/Y _08308_/A _08441_/X VGND VGND VPWR VPWR _08697_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_90_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08392_ _08392_/A VGND VGND VPWR VPWR _08392_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09013_ _08893_/X _09021_/S _08579_/Y VGND VGND VPWR VPWR _09020_/S sky130_fd_sc_hd__o21ai_1
XFILLER_117_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09915_ _09859_/A _09859_/B _09914_/Y VGND VGND VPWR VPWR _10946_/A sky130_fd_sc_hd__a21oi_1
XFILLER_86_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09846_ _10491_/B _10490_/A VGND VGND VPWR VPWR _09846_/X sky130_fd_sc_hd__or2_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09777_ _10079_/A _09775_/Y _09776_/Y VGND VGND VPWR VPWR _09779_/B sky130_fd_sc_hd__o21ai_2
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08728_ _08715_/A _08715_/B _08715_/X _08727_/X VGND VGND VPWR VPWR _08729_/A sky130_fd_sc_hd__a22o_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _10099_/B VGND VGND VPWR VPWR _08679_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11573_/Y _11669_/X _11573_/Y _11669_/X VGND VGND VPWR VPWR _11673_/B sky130_fd_sc_hd__a2bb2o_1
X_10621_ _12232_/A _11792_/B VGND VGND VPWR VPWR _12916_/A sky130_fd_sc_hd__or2_1
XFILLER_10_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13340_ _13340_/A _13340_/B VGND VGND VPWR VPWR _13340_/X sky130_fd_sc_hd__and2_1
X_10552_ _10552_/A _11810_/A VGND VGND VPWR VPWR _10552_/Y sky130_fd_sc_hd__nor2_1
X_13271_ _12043_/A _13270_/Y _12043_/A _13270_/Y VGND VGND VPWR VPWR _13272_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12222_ _12222_/A _12141_/X VGND VGND VPWR VPWR _12222_/X sky130_fd_sc_hd__or2b_1
X_15010_ _15044_/A _15044_/B VGND VGND VPWR VPWR _15058_/A sky130_fd_sc_hd__and2_1
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10483_ _09848_/A _09848_/B _09851_/A VGND VGND VPWR VPWR _10483_/X sky130_fd_sc_hd__o21ba_1
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12153_ _13898_/A _12153_/B VGND VGND VPWR VPWR _12153_/X sky130_fd_sc_hd__or2_1
XFILLER_96_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12084_ _12084_/A VGND VGND VPWR VPWR _12174_/B sky130_fd_sc_hd__inv_2
X_11104_ _09782_/A _09380_/A _09432_/X VGND VGND VPWR VPWR _11105_/A sky130_fd_sc_hd__o21ai_1
X_15912_ _15978_/A _15978_/B VGND VGND VPWR VPWR _15912_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11035_ _13560_/A VGND VGND VPWR VPWR _12844_/A sky130_fd_sc_hd__buf_1
X_15843_ _14220_/A _15842_/X _12621_/X VGND VGND VPWR VPWR _15843_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15774_ _15774_/A _16028_/A VGND VGND VPWR VPWR _15774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12986_ _13693_/A VGND VGND VPWR VPWR _14489_/A sky130_fd_sc_hd__inv_2
XFILLER_64_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14725_ _14725_/A _14725_/B VGND VGND VPWR VPWR _14807_/B sky130_fd_sc_hd__and2_1
X_11937_ _13699_/A _11978_/B _11936_/Y VGND VGND VPWR VPWR _11937_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14656_ _15341_/A _14656_/B VGND VGND VPWR VPWR _14656_/Y sky130_fd_sc_hd__nand2_1
X_11868_ _13633_/A _11909_/B _11867_/Y VGND VGND VPWR VPWR _11868_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14587_ _14543_/Y _14585_/X _14586_/Y VGND VGND VPWR VPWR _14587_/X sky130_fd_sc_hd__o21a_1
X_13607_ _13607_/A _13574_/X VGND VGND VPWR VPWR _13607_/X sky130_fd_sc_hd__or2b_1
X_11799_ _11799_/A VGND VGND VPWR VPWR _11799_/Y sky130_fd_sc_hd__inv_2
X_10819_ _10819_/A VGND VGND VPWR VPWR _10819_/Y sky130_fd_sc_hd__inv_2
X_16326_ _16326_/A _16326_/B VGND VGND VPWR VPWR _16326_/Y sky130_fd_sc_hd__nand2_1
X_13538_ _15040_/A _13513_/B _13513_/Y _13537_/X VGND VGND VPWR VPWR _13538_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16257_ _16257_/A VGND VGND VPWR VPWR _16324_/A sky130_fd_sc_hd__buf_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13469_ _13467_/Y _13468_/X _13467_/Y _13468_/X VGND VGND VPWR VPWR _13469_/X sky130_fd_sc_hd__a2bb2o_1
X_16188_ _16105_/X _16187_/X _16105_/X _16187_/X VGND VGND VPWR VPWR _16189_/B sky130_fd_sc_hd__a2bb2oi_1
X_15208_ _15208_/A _15208_/B VGND VGND VPWR VPWR _15208_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15139_ _15089_/X _15138_/Y _15089_/X _15138_/Y VGND VGND VPWR VPWR _15140_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09700_ _09700_/A VGND VGND VPWR VPWR _09700_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09631_ _09952_/A _09631_/B VGND VGND VPWR VPWR _09632_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09562_ _09567_/A _09560_/X _09567_/B VGND VGND VPWR VPWR _09562_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_82_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08513_ _09863_/A _08509_/A _08464_/A _08512_/X _08464_/Y VGND VGND VPWR VPWR _08989_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_70_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09493_ _08806_/A _09466_/X _08806_/A _09466_/X VGND VGND VPWR VPWR _09494_/B sky130_fd_sc_hd__o2bb2a_1
X_08444_ _08711_/A VGND VGND VPWR VPWR _09333_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08375_ input4/X _08248_/B _08317_/B _08447_/A VGND VGND VPWR VPWR _08454_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09829_ _09829_/A _09829_/B VGND VGND VPWR VPWR _09830_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12840_ _12840_/A _12840_/B VGND VGND VPWR VPWR _12840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12771_/A _12771_/B VGND VGND VPWR VPWR _12771_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15490_ _15485_/X _15489_/X _15485_/X _15489_/X VGND VGND VPWR VPWR _15552_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _15211_/A _14510_/B VGND VGND VPWR VPWR _14510_/X sky130_fd_sc_hd__or2_1
X_11722_ _10282_/A _11721_/Y _10899_/B _10347_/A VGND VGND VPWR VPWR _11733_/B sky130_fd_sc_hd__o22a_1
XFILLER_30_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11653_/A VGND VGND VPWR VPWR _13989_/A sky130_fd_sc_hd__buf_1
X_14441_ _14436_/X _14440_/X _14436_/X _14440_/X VGND VGND VPWR VPWR _14469_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14372_ _14372_/A _14372_/B VGND VGND VPWR VPWR _14373_/A sky130_fd_sc_hd__or2_1
XFILLER_80_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10604_ _11837_/A _10527_/B _10527_/Y VGND VGND VPWR VPWR _10604_/Y sky130_fd_sc_hd__o21ai_1
X_16111_ _16073_/X _16109_/X _16171_/B VGND VGND VPWR VPWR _16111_/X sky130_fd_sc_hd__o21a_1
X_13323_ _14737_/A _13294_/B _13294_/Y VGND VGND VPWR VPWR _13323_/Y sky130_fd_sc_hd__o21ai_1
X_11584_ _13139_/A VGND VGND VPWR VPWR _11653_/A sky130_fd_sc_hd__inv_2
X_10535_ _09898_/A _09898_/B _09901_/A VGND VGND VPWR VPWR _10535_/X sky130_fd_sc_hd__o21ba_1
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16042_ _16042_/A _16042_/B VGND VGND VPWR VPWR _16042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13254_ _13189_/X _13253_/Y _13189_/X _13253_/Y VGND VGND VPWR VPWR _13282_/B sky130_fd_sc_hd__a2bb2o_1
X_10466_ _11854_/A _10554_/B _10465_/Y VGND VGND VPWR VPWR _10467_/A sky130_fd_sc_hd__o21ai_2
XFILLER_108_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12205_ _12152_/X _12204_/X _12152_/X _12204_/X VGND VGND VPWR VPWR _12206_/B sky130_fd_sc_hd__a2bb2o_1
X_13185_ _13178_/Y _13183_/X _13184_/Y VGND VGND VPWR VPWR _13185_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12136_ _13936_/A _13936_/B _12134_/X _12233_/A VGND VGND VPWR VPWR _12136_/X sky130_fd_sc_hd__a31o_1
XFILLER_69_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10397_ _11775_/A VGND VGND VPWR VPWR _13564_/A sky130_fd_sc_hd__buf_1
XFILLER_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12067_ _12066_/Y _11977_/X _12011_/Y VGND VGND VPWR VPWR _12067_/X sky130_fd_sc_hd__o21a_1
X_11018_ _11018_/A _10919_/X VGND VGND VPWR VPWR _11018_/X sky130_fd_sc_hd__or2b_1
XFILLER_65_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15826_ _15697_/X _15825_/Y _15703_/Y VGND VGND VPWR VPWR _15826_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15757_ _14911_/X _15756_/X _14911_/X _15756_/X VGND VGND VPWR VPWR _15758_/B sky130_fd_sc_hd__a2bb2oi_1
X_12969_ _14592_/A _13028_/B VGND VGND VPWR VPWR _13055_/A sky130_fd_sc_hd__and2_1
XFILLER_18_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15688_ _14400_/Y _15687_/X _14400_/Y _15687_/X VGND VGND VPWR VPWR _15694_/B sky130_fd_sc_hd__a2bb2o_1
X_14708_ _14729_/A _14729_/B VGND VGND VPWR VPWR _14800_/A sky130_fd_sc_hd__and2_1
X_14639_ _15272_/A _14574_/B _14574_/Y VGND VGND VPWR VPWR _14639_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16309_ _16251_/A _16309_/A2 _16251_/Y VGND VGND VPWR VPWR _16309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08993_ _09341_/A _08748_/Y _09342_/A VGND VGND VPWR VPWR _08993_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09614_ _09548_/X _09613_/Y _09548_/X _09613_/Y VGND VGND VPWR VPWR _09652_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09545_ _09538_/A _09538_/B _09538_/X _09544_/X VGND VGND VPWR VPWR _09546_/A sky130_fd_sc_hd__o22a_1
X_09476_ _10009_/A _09476_/B VGND VGND VPWR VPWR _09476_/X sky130_fd_sc_hd__or2_1
X_08427_ _08714_/A VGND VGND VPWR VPWR _08794_/A sky130_fd_sc_hd__buf_1
XFILLER_12_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08358_ _08358_/A input18/X VGND VGND VPWR VPWR _08399_/A sky130_fd_sc_hd__nor2_1
X_08289_ _08336_/A input31/X _08337_/A _08339_/A VGND VGND VPWR VPWR _08334_/A sky130_fd_sc_hd__o22a_1
XFILLER_118_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10320_ _09958_/A _09958_/B _09958_/Y VGND VGND VPWR VPWR _10320_/Y sky130_fd_sc_hd__o21ai_1
X_10251_ _10251_/A VGND VGND VPWR VPWR _10251_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10182_ _10182_/A VGND VGND VPWR VPWR _10182_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14990_ _12430_/X _14989_/X _12430_/X _14989_/X VGND VGND VPWR VPWR _14990_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_115_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13941_ _14041_/A _13939_/X _13940_/X VGND VGND VPWR VPWR _13941_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13872_ _13872_/A _13873_/B VGND VGND VPWR VPWR _13874_/A sky130_fd_sc_hd__and2_1
XFILLER_47_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15611_ _16040_/A VGND VGND VPWR VPWR _15677_/A sky130_fd_sc_hd__inv_2
XFILLER_62_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12823_ _12763_/A _12763_/B _12763_/Y VGND VGND VPWR VPWR _12823_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15542_ _15542_/A _15542_/B VGND VGND VPWR VPWR _15542_/X sky130_fd_sc_hd__or2_1
XFILLER_91_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12754_ _12703_/A _12703_/B _12703_/A _12703_/B VGND VGND VPWR VPWR _12754_/X sky130_fd_sc_hd__a2bb2o_1
X_11705_ _11705_/A VGND VGND VPWR VPWR _11706_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15473_ _15473_/A _15473_/B VGND VGND VPWR VPWR _15473_/Y sky130_fd_sc_hd__nand2_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _11152_/A _12672_/A _11152_/Y _12672_/Y VGND VGND VPWR VPWR _12686_/B sky130_fd_sc_hd__o22a_1
X_11636_ _12863_/A _11636_/B VGND VGND VPWR VPWR _11636_/X sky130_fd_sc_hd__or2_1
X_14424_ _11773_/Y _14417_/X _11773_/Y _14417_/X VGND VGND VPWR VPWR _14425_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14355_ _15881_/A _14251_/B _14251_/Y VGND VGND VPWR VPWR _14355_/Y sky130_fd_sc_hd__o21ai_1
X_11567_ _08986_/A _08986_/B _08986_/Y VGND VGND VPWR VPWR _11567_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14286_ _14286_/A _15908_/A VGND VGND VPWR VPWR _14286_/X sky130_fd_sc_hd__or2_1
X_13306_ _14858_/A _13306_/B VGND VGND VPWR VPWR _13306_/Y sky130_fd_sc_hd__nand2_1
X_10518_ _11791_/A _10430_/B _11791_/A _10430_/B VGND VGND VPWR VPWR _10518_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16025_ _16030_/A _16030_/B VGND VGND VPWR VPWR _16025_/Y sky130_fd_sc_hd__nor2_1
X_13237_ _14474_/A VGND VGND VPWR VPWR _14735_/A sky130_fd_sc_hd__buf_1
X_11498_ _12365_/A _11498_/B VGND VGND VPWR VPWR _11498_/Y sky130_fd_sc_hd__nor2_1
X_10449_ _10451_/A VGND VGND VPWR VPWR _10449_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13168_ _13190_/A _13190_/B VGND VGND VPWR VPWR _13168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12119_ _13914_/A _12145_/B VGND VGND VPWR VPWR _12216_/A sky130_fd_sc_hd__and2_1
X_13099_ _13007_/A _13098_/Y _13007_/A _13098_/Y VGND VGND VPWR VPWR _13101_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15809_ _16108_/A _15809_/B VGND VGND VPWR VPWR _15809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09330_ _09330_/A _09330_/B VGND VGND VPWR VPWR _09330_/Y sky130_fd_sc_hd__nand2_1
X_09261_ _09260_/X _08894_/Y _09260_/X _08894_/Y VGND VGND VPWR VPWR _10242_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09192_ _09561_/B _09156_/X _09190_/Y _11664_/B VGND VGND VPWR VPWR _09193_/A sky130_fd_sc_hd__o22a_1
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08976_ _08976_/A _08976_/B VGND VGND VPWR VPWR _11371_/B sky130_fd_sc_hd__or2_1
XFILLER_75_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09528_ _09528_/A VGND VGND VPWR VPWR _09528_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09459_ _09459_/A _09459_/B VGND VGND VPWR VPWR _09459_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12470_ _13973_/A _12447_/B _12447_/Y _12450_/X VGND VGND VPWR VPWR _12470_/Y sky130_fd_sc_hd__o2bb2ai_1
X_11421_ _13406_/A _13406_/B _12606_/B _11420_/X VGND VGND VPWR VPWR _11422_/B sky130_fd_sc_hd__a31o_1
X_14140_ _14134_/X _14137_/Y _14864_/A _14139_/Y VGND VGND VPWR VPWR _14140_/X sky130_fd_sc_hd__o22a_1
X_11352_ _11267_/X _11351_/X _11267_/X _11351_/X VGND VGND VPWR VPWR _11353_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10303_ _10303_/A VGND VGND VPWR VPWR _11759_/A sky130_fd_sc_hd__inv_2
XFILLER_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14071_ _14956_/A _13989_/B _13989_/Y _13992_/X VGND VGND VPWR VPWR _14071_/X sky130_fd_sc_hd__o2bb2a_1
X_11283_ _13048_/A _11170_/B _11170_/Y _11110_/X VGND VGND VPWR VPWR _11283_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13022_ _14481_/A _13022_/B VGND VGND VPWR VPWR _13022_/X sky130_fd_sc_hd__or2_1
X_10234_ _10234_/A VGND VGND VPWR VPWR _10234_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10165_ _10167_/A VGND VGND VPWR VPWR _10469_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14973_ _12428_/A _12421_/Y _12432_/Y _14936_/X VGND VGND VPWR VPWR _14973_/Y sky130_fd_sc_hd__o22ai_2
X_10096_ _10215_/A _11237_/A VGND VGND VPWR VPWR _11733_/A sky130_fd_sc_hd__or2_1
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13924_ _13843_/X _13923_/Y _13843_/X _13923_/Y VGND VGND VPWR VPWR _13944_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13855_ _13809_/Y _13853_/X _13854_/Y VGND VGND VPWR VPWR _13855_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12806_ _12774_/X _12805_/Y _12774_/X _12805_/Y VGND VGND VPWR VPWR _12850_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10998_ _13053_/A _10998_/B VGND VGND VPWR VPWR _10998_/Y sky130_fd_sc_hd__nand2_1
X_13786_ _13786_/A _13786_/B VGND VGND VPWR VPWR _13868_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15525_ _15521_/Y _15632_/A _15524_/Y VGND VGND VPWR VPWR _15529_/B sky130_fd_sc_hd__o21ai_2
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12715_/X _12736_/X _12715_/X _12736_/X VGND VGND VPWR VPWR _12777_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15456_ _15456_/A _15406_/X VGND VGND VPWR VPWR _15456_/X sky130_fd_sc_hd__or2b_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _12668_/A VGND VGND VPWR VPWR _12668_/Y sky130_fd_sc_hd__inv_2
X_14407_ _12651_/Y _14406_/X _12651_/Y _14406_/X VGND VGND VPWR VPWR _14407_/Y sky130_fd_sc_hd__a2bb2oi_1
X_11619_ _12416_/A VGND VGND VPWR VPWR _12379_/A sky130_fd_sc_hd__inv_2
XFILLER_129_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12599_ _12594_/Y _12598_/A _12594_/A _12598_/Y _11705_/A VGND VGND VPWR VPWR _12617_/A
+ sky130_fd_sc_hd__o221a_1
X_15387_ _15387_/A _15333_/X VGND VGND VPWR VPWR _15387_/X sky130_fd_sc_hd__or2b_1
X_14338_ _14259_/A _14337_/Y _14259_/A _14337_/Y VGND VGND VPWR VPWR _14384_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14269_ _15863_/A _14269_/B VGND VGND VPWR VPWR _14269_/Y sky130_fd_sc_hd__nand2_1
X_16008_ _16008_/A _15958_/X VGND VGND VPWR VPWR _16008_/X sky130_fd_sc_hd__or2b_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08830_/A VGND VGND VPWR VPWR _08831_/A sky130_fd_sc_hd__inv_2
XFILLER_112_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08761_ _10009_/A VGND VGND VPWR VPWR _08762_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08692_ _08692_/A _10119_/B VGND VGND VPWR VPWR _08876_/B sky130_fd_sc_hd__and2_1
XFILLER_81_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09313_ _09313_/A _09313_/B VGND VGND VPWR VPWR _09313_/Y sky130_fd_sc_hd__nand2_1
X_09244_ _09467_/B _09857_/A _09212_/Y _09243_/X VGND VGND VPWR VPWR _09244_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09175_ _09432_/A _09175_/B VGND VGND VPWR VPWR _09175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08959_ _08681_/Y _08958_/X _08681_/Y _08958_/X VGND VGND VPWR VPWR _11397_/A sky130_fd_sc_hd__o2bb2a_1
X_11970_ _11970_/A _11970_/B VGND VGND VPWR VPWR _11970_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10921_ _10921_/A VGND VGND VPWR VPWR _14611_/A sky130_fd_sc_hd__buf_1
XFILLER_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10852_ _10918_/A _10919_/B VGND VGND VPWR VPWR _11018_/A sky130_fd_sc_hd__and2_1
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13640_ _13640_/A VGND VGND VPWR VPWR _13640_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10783_ _10781_/Y _10782_/Y _10701_/Y VGND VGND VPWR VPWR _10936_/A sky130_fd_sc_hd__o21ai_1
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _13531_/X _13570_/Y _13531_/X _13570_/Y VGND VGND VPWR VPWR _13574_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16290_ _16332_/A _16332_/B VGND VGND VPWR VPWR _16290_/Y sky130_fd_sc_hd__nor2_1
X_12522_ _12522_/A _12522_/B VGND VGND VPWR VPWR _12522_/Y sky130_fd_sc_hd__nand2_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15310_ _15277_/X _15309_/Y _15277_/X _15309_/Y VGND VGND VPWR VPWR _15341_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15241_ _15187_/A _15187_/B _15187_/Y VGND VGND VPWR VPWR _15241_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12453_ _13979_/A _12452_/B _12452_/Y VGND VGND VPWR VPWR _12453_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11404_ _12329_/A VGND VGND VPWR VPWR _15519_/A sky130_fd_sc_hd__buf_1
X_15172_ _15171_/A _15425_/B _15171_/Y VGND VGND VPWR VPWR _15172_/Y sky130_fd_sc_hd__o21ai_1
X_12384_ _12435_/B _12383_/Y _12435_/B _12383_/Y VGND VGND VPWR VPWR _12440_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14123_ _14123_/A _14060_/X VGND VGND VPWR VPWR _14123_/X sky130_fd_sc_hd__or2b_1
X_11335_ _11305_/X _11334_/X _11305_/X _11334_/X VGND VGND VPWR VPWR _11504_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14054_ _15458_/A _14028_/B _14028_/X _14053_/X VGND VGND VPWR VPWR _14054_/X sky130_fd_sc_hd__o22a_1
X_11266_ _14009_/A VGND VGND VPWR VPWR _14064_/A sky130_fd_sc_hd__buf_1
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13005_ _13002_/X _13004_/X _13002_/X _13004_/X VGND VGND VPWR VPWR _13008_/B sky130_fd_sc_hd__a2bb2o_1
X_10217_ _10059_/A _10059_/B _10059_/Y VGND VGND VPWR VPWR _10217_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11197_ _14058_/A _11197_/B VGND VGND VPWR VPWR _11197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10148_ _10117_/A _10117_/B _10118_/A VGND VGND VPWR VPWR _10151_/A sky130_fd_sc_hd__a21bo_1
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14956_ _14956_/A _14956_/B VGND VGND VPWR VPWR _14956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10079_ _10079_/A _10079_/B VGND VGND VPWR VPWR _10813_/B sky130_fd_sc_hd__or2_1
X_13907_ _14615_/A _13852_/B _13852_/Y VGND VGND VPWR VPWR _13907_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14887_ _14798_/A _14798_/B _14798_/A _14798_/B VGND VGND VPWR VPWR _14887_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13838_ _13838_/A _13838_/B VGND VGND VPWR VPWR _13838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13769_ _13769_/A _13769_/B VGND VGND VPWR VPWR _13769_/X sky130_fd_sc_hd__or2_1
X_15508_ _12235_/X _15507_/Y _12235_/X _15507_/Y VGND VGND VPWR VPWR _15509_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15439_ _15417_/X _15438_/X _15417_/X _15438_/X VGND VGND VPWR VPWR _15440_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09931_ _09931_/A _09930_/Y VGND VGND VPWR VPWR _09932_/B sky130_fd_sc_hd__or2b_1
XFILLER_131_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09862_ _09862_/A _09924_/A VGND VGND VPWR VPWR _09863_/B sky130_fd_sc_hd__or2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08813_ _08813_/A VGND VGND VPWR VPWR _08814_/A sky130_fd_sc_hd__inv_2
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09793_/A _09793_/B VGND VGND VPWR VPWR _09794_/A sky130_fd_sc_hd__or2_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08744_ _08709_/Y _08742_/Y _08743_/X VGND VGND VPWR VPWR _08745_/A sky130_fd_sc_hd__o21ai_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08675_ _08664_/X _08402_/X _10228_/A _08674_/Y VGND VGND VPWR VPWR _10098_/B sky130_fd_sc_hd__a31o_1
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09227_ _09458_/B _09690_/A VGND VGND VPWR VPWR _09227_/X sky130_fd_sc_hd__or2_1
X_09158_ _09158_/A VGND VGND VPWR VPWR _09158_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09089_ _10015_/B _09074_/B _09075_/B VGND VGND VPWR VPWR _09701_/A sky130_fd_sc_hd__a21bo_1
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11120_ _09966_/Y _11119_/A _10083_/A _11119_/Y _11590_/A VGND VGND VPWR VPWR _12254_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11051_ _10910_/X _11050_/X _10910_/X _11050_/X VGND VGND VPWR VPWR _11079_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10002_ _09521_/Y _09792_/A _09521_/Y _09792_/A VGND VGND VPWR VPWR _10002_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14810_ _15398_/A _14718_/B _15398_/A _14718_/B VGND VGND VPWR VPWR _14810_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15790_ _15793_/A _15794_/B VGND VGND VPWR VPWR _15790_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14741_ _14741_/A _14741_/B VGND VGND VPWR VPWR _14741_/X sky130_fd_sc_hd__or2_1
X_11953_ _11894_/A _11952_/Y _11894_/A _11952_/Y VGND VGND VPWR VPWR _11966_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10904_ _10904_/A _11411_/A VGND VGND VPWR VPWR _12041_/B sky130_fd_sc_hd__or2_1
XFILLER_72_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11884_ _11834_/X _11883_/Y _11834_/X _11883_/Y VGND VGND VPWR VPWR _11892_/B sky130_fd_sc_hd__a2bb2o_1
X_14672_ _15044_/A _12168_/Y _12090_/Y _14595_/X VGND VGND VPWR VPWR _14672_/X sky130_fd_sc_hd__o22a_1
XFILLER_45_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16411_ _16454_/A _16411_/B VGND VGND VPWR VPWR _16474_/D sky130_fd_sc_hd__or2_1
X_13623_ _13602_/Y _13620_/X _13622_/Y VGND VGND VPWR VPWR _13624_/A sky130_fd_sc_hd__o21ai_2
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10835_ _10796_/X _10834_/X _10796_/X _10834_/X VGND VGND VPWR VPWR _10944_/B sky130_fd_sc_hd__a2bb2o_1
X_16342_ _16361_/A VGND VGND VPWR VPWR _16343_/A sky130_fd_sc_hd__buf_1
X_10766_ _11958_/A _10766_/B VGND VGND VPWR VPWR _10766_/X sky130_fd_sc_hd__or2_1
X_13554_ _15036_/A _13519_/B _13519_/Y VGND VGND VPWR VPWR _13554_/Y sky130_fd_sc_hd__o21ai_1
X_16273_ _16273_/A _16338_/A VGND VGND VPWR VPWR _16273_/Y sky130_fd_sc_hd__nand2_1
X_12505_ _13446_/A _11356_/B _11356_/Y VGND VGND VPWR VPWR _12506_/B sky130_fd_sc_hd__o21a_1
X_10697_ _10658_/X _10696_/X _10658_/X _10696_/X VGND VGND VPWR VPWR _10789_/B sky130_fd_sc_hd__a2bb2o_1
X_13485_ _10449_/Y _11764_/A _10387_/Y _13484_/X VGND VGND VPWR VPWR _13485_/X sky130_fd_sc_hd__o22a_1
XFILLER_126_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15224_ _15193_/A _15193_/B _15193_/Y _15223_/X VGND VGND VPWR VPWR _15224_/X sky130_fd_sc_hd__a2bb2o_1
X_12436_ _12785_/A _12435_/B _12435_/Y _12382_/B VGND VGND VPWR VPWR _12437_/B sky130_fd_sc_hd__a2bb2o_1
X_15155_ _15122_/A _15122_/B _15122_/Y _15154_/X VGND VGND VPWR VPWR _15155_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14106_ _14106_/A _14106_/B VGND VGND VPWR VPWR _14106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12367_ _13786_/A _12367_/B VGND VGND VPWR VPWR _12367_/X sky130_fd_sc_hd__and2_1
X_12298_ _14009_/A _12297_/B _12297_/Y VGND VGND VPWR VPWR _12298_/Y sky130_fd_sc_hd__o21ai_1
X_15086_ _15087_/A _15087_/B VGND VGND VPWR VPWR _15144_/A sky130_fd_sc_hd__and2_1
X_11318_ _11604_/A _11318_/B VGND VGND VPWR VPWR _11319_/A sky130_fd_sc_hd__or2_1
X_11249_ _11411_/A _11249_/B _13936_/B VGND VGND VPWR VPWR _11249_/X sky130_fd_sc_hd__or3_1
X_14037_ _15400_/A _13942_/B _13942_/Y VGND VGND VPWR VPWR _14037_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15988_ _15988_/A _15982_/X VGND VGND VPWR VPWR _15988_/X sky130_fd_sc_hd__or2b_1
XFILLER_48_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14939_ _14934_/A _14938_/B _14938_/Y VGND VGND VPWR VPWR _14939_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08460_ _08460_/A VGND VGND VPWR VPWR _08460_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08391_ input9/X _08279_/B _08279_/Y VGND VGND VPWR VPWR _08392_/A sky130_fd_sc_hd__a21oi_2
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09012_ _08795_/X _09011_/Y _09213_/B VGND VGND VPWR VPWR _09021_/S sky130_fd_sc_hd__a21oi_1
XFILLER_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09914_ _09914_/A VGND VGND VPWR VPWR _09914_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09845_ _09801_/A _09801_/B _09844_/Y VGND VGND VPWR VPWR _10490_/A sky130_fd_sc_hd__a21oi_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09776_ _09776_/A _09776_/B VGND VGND VPWR VPWR _09776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08727_ _08716_/A _08716_/B _08716_/X _08726_/X VGND VGND VPWR VPWR _08727_/X sky130_fd_sc_hd__a22o_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08658_ _08657_/Y _08403_/Y _08657_/Y _08403_/Y VGND VGND VPWR VPWR _10099_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08589_ _08589_/A _08589_/B VGND VGND VPWR VPWR _09455_/B sky130_fd_sc_hd__or2_1
X_10620_ _10620_/A _10622_/C VGND VGND VPWR VPWR _10623_/A sky130_fd_sc_hd__nor2_1
X_10551_ _11852_/A VGND VGND VPWR VPWR _11810_/A sky130_fd_sc_hd__inv_2
X_13270_ _15329_/A _13182_/B _13182_/Y VGND VGND VPWR VPWR _13270_/Y sky130_fd_sc_hd__a21oi_1
X_10482_ _13629_/A _10533_/B VGND VGND VPWR VPWR _10482_/Y sky130_fd_sc_hd__nor2_1
X_12221_ _12221_/A _12221_/B VGND VGND VPWR VPWR _12221_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12152_ _12207_/A _12150_/X _12151_/X VGND VGND VPWR VPWR _12152_/X sky130_fd_sc_hd__o21a_1
X_11103_ _11004_/A _10923_/X _11003_/X VGND VGND VPWR VPWR _11103_/X sky130_fd_sc_hd__o21a_1
XFILLER_78_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12083_ _10816_/A _11994_/A _10964_/B _12082_/Y VGND VGND VPWR VPWR _12084_/A sky130_fd_sc_hd__o22a_1
X_15911_ _14171_/X _15851_/X _14171_/X _15851_/X VGND VGND VPWR VPWR _15978_/B sky130_fd_sc_hd__a2bb2o_1
X_11034_ _13914_/A _11085_/B VGND VGND VPWR VPWR _11216_/A sky130_fd_sc_hd__and2_1
XFILLER_78_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15842_ _14226_/A _15841_/X _12619_/X VGND VGND VPWR VPWR _15842_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15773_ _16084_/A VGND VGND VPWR VPWR _15782_/A sky130_fd_sc_hd__inv_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12985_ _14485_/A _13020_/B VGND VGND VPWR VPWR _13075_/A sky130_fd_sc_hd__and2_1
XFILLER_45_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14724_ _15398_/A _14718_/B _14718_/X _14723_/X VGND VGND VPWR VPWR _14724_/X sky130_fd_sc_hd__o22a_1
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11936_ _11978_/A _11978_/B VGND VGND VPWR VPWR _11936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14655_ _14626_/Y _14653_/X _14654_/Y VGND VGND VPWR VPWR _14655_/X sky130_fd_sc_hd__o21a_1
X_11867_ _11867_/A _11909_/B VGND VGND VPWR VPWR _11867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14586_ _14586_/A _14586_/B VGND VGND VPWR VPWR _14586_/Y sky130_fd_sc_hd__nand2_1
X_13606_ _13606_/A _13606_/B VGND VGND VPWR VPWR _13606_/Y sky130_fd_sc_hd__nor2_1
X_11798_ _11798_/A _11798_/B VGND VGND VPWR VPWR _11798_/X sky130_fd_sc_hd__or2_1
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10818_ _10818_/A VGND VGND VPWR VPWR _10818_/Y sky130_fd_sc_hd__inv_2
X_16325_ _16302_/Y _16323_/X _16324_/Y VGND VGND VPWR VPWR _16325_/X sky130_fd_sc_hd__o21a_1
X_13537_ _15038_/A _13516_/B _13516_/Y _13536_/X VGND VGND VPWR VPWR _13537_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10749_ _10749_/A VGND VGND VPWR VPWR _10749_/Y sky130_fd_sc_hd__inv_2
X_16256_ _16211_/Y _16254_/X _16255_/Y VGND VGND VPWR VPWR _16256_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13468_ _15289_/A _13139_/B _13139_/Y _13207_/X VGND VGND VPWR VPWR _13468_/X sky130_fd_sc_hd__o2bb2a_1
X_15207_ _15148_/X _15206_/Y _15148_/X _15206_/Y VGND VGND VPWR VPWR _15208_/B sky130_fd_sc_hd__a2bb2o_1
X_16187_ _16079_/X _16187_/B VGND VGND VPWR VPWR _16187_/X sky130_fd_sc_hd__and2b_1
X_13399_ _14093_/A VGND VGND VPWR VPWR _14096_/A sky130_fd_sc_hd__buf_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12419_ _12419_/A _12419_/B VGND VGND VPWR VPWR _12419_/Y sky130_fd_sc_hd__nand2_1
X_15138_ _15081_/A _15081_/B _15081_/Y VGND VGND VPWR VPWR _15138_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15069_ _15069_/A _15069_/B VGND VGND VPWR VPWR _15069_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09630_ _09707_/A _09628_/Y _08929_/B _09629_/X VGND VGND VPWR VPWR _09631_/B sky130_fd_sc_hd__o22a_1
XFILLER_83_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09561_ _09561_/A _09561_/B VGND VGND VPWR VPWR _09567_/B sky130_fd_sc_hd__and2_1
XFILLER_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08512_ _09346_/B _09791_/C VGND VGND VPWR VPWR _08512_/X sky130_fd_sc_hd__or2_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09492_ _09492_/A _09492_/B VGND VGND VPWR VPWR _09492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08443_ _08554_/A VGND VGND VPWR VPWR _08711_/A sky130_fd_sc_hd__inv_2
X_08374_ input3/X _08251_/B _08322_/B _08440_/A VGND VGND VPWR VPWR _08447_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09828_ _10102_/A _09829_/A _09503_/B _09827_/X VGND VGND VPWR VPWR _09832_/A sky130_fd_sc_hd__a31o_1
XFILLER_73_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09759_ _10043_/A VGND VGND VPWR VPWR _10083_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12750_/Y _12768_/X _12769_/Y VGND VGND VPWR VPWR _12770_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11721_/A _11721_/B VGND VGND VPWR VPWR _11721_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11653_/A _11654_/B VGND VGND VPWR VPWR _11655_/A sky130_fd_sc_hd__and2_1
X_14440_ _14439_/A _14439_/B _14439_/Y VGND VGND VPWR VPWR _14440_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14371_ _15838_/A VGND VGND VPWR VPWR _14371_/X sky130_fd_sc_hd__buf_1
X_10603_ _09951_/Y _10602_/Y _10216_/X _10602_/A _09797_/A VGND VGND VPWR VPWR _10744_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16110_ _16110_/A _16110_/B VGND VGND VPWR VPWR _16171_/B sky130_fd_sc_hd__or2_1
X_13322_ _13367_/A _13367_/B VGND VGND VPWR VPWR _13385_/A sky130_fd_sc_hd__and2_1
X_11583_ _11583_/A _11583_/B VGND VGND VPWR VPWR _13139_/A sky130_fd_sc_hd__or2_2
X_10534_ _10482_/Y _10532_/X _10533_/Y VGND VGND VPWR VPWR _10534_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16041_ _16010_/Y _16039_/X _16040_/Y VGND VGND VPWR VPWR _16041_/X sky130_fd_sc_hd__o21a_1
X_13253_ _13190_/A _13190_/B _13190_/Y VGND VGND VPWR VPWR _13253_/Y sky130_fd_sc_hd__o21ai_1
X_10465_ _11854_/A _10554_/B VGND VGND VPWR VPWR _10465_/Y sky130_fd_sc_hd__nand2_1
X_12204_ _12204_/A _12153_/X VGND VGND VPWR VPWR _12204_/X sky130_fd_sc_hd__or2b_1
X_13184_ _13829_/A _13184_/B VGND VGND VPWR VPWR _13184_/Y sky130_fd_sc_hd__nand2_1
X_10396_ _10396_/A VGND VGND VPWR VPWR _11775_/A sky130_fd_sc_hd__buf_1
XFILLER_97_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12135_ _12135_/A _12135_/B VGND VGND VPWR VPWR _12233_/A sky130_fd_sc_hd__and2_1
XFILLER_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12066_ _12066_/A _12066_/B VGND VGND VPWR VPWR _12066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11017_ _15066_/A VGND VGND VPWR VPWR _13906_/A sky130_fd_sc_hd__buf_1
XFILLER_77_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15825_ _15991_/A _15825_/B VGND VGND VPWR VPWR _15825_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15756_ _14912_/A _14912_/B _14912_/Y VGND VGND VPWR VPWR _15756_/X sky130_fd_sc_hd__o21a_1
X_12968_ _12939_/X _12967_/Y _12939_/X _12967_/Y VGND VGND VPWR VPWR _13028_/B sky130_fd_sc_hd__a2bb2o_1
X_15687_ _15687_/A _14401_/X VGND VGND VPWR VPWR _15687_/X sky130_fd_sc_hd__or2b_1
X_14707_ _14651_/X _14706_/Y _14651_/X _14706_/Y VGND VGND VPWR VPWR _14729_/B sky130_fd_sc_hd__a2bb2o_1
X_12899_ _14465_/A _12930_/B VGND VGND VPWR VPWR _12899_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11919_ _11918_/A _11918_/B _11918_/X _11859_/B VGND VGND VPWR VPWR _11990_/B sky130_fd_sc_hd__a22o_1
X_14638_ _15333_/A _14648_/B VGND VGND VPWR VPWR _14638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16308_ _16320_/A _16320_/B VGND VGND VPWR VPWR _16308_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14569_ _15216_/A _14508_/B _14508_/Y VGND VGND VPWR VPWR _14569_/Y sky130_fd_sc_hd__a21oi_1
X_16239_ _16249_/B VGND VGND VPWR VPWR _16240_/B sky130_fd_sc_hd__buf_1
X_08992_ _09518_/A _10134_/A _08752_/X _08868_/Y VGND VGND VPWR VPWR _08992_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09613_ _09613_/A _09613_/B VGND VGND VPWR VPWR _09613_/Y sky130_fd_sc_hd__nor2_1
X_09544_ _09539_/A _09539_/B _09539_/X _09543_/X VGND VGND VPWR VPWR _09544_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09475_ _09450_/Y _09473_/X _09474_/X VGND VGND VPWR VPWR _09475_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08426_ _09213_/A VGND VGND VPWR VPWR _08714_/A sky130_fd_sc_hd__inv_2
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08357_ input26/X _08357_/B VGND VGND VPWR VPWR _08387_/B sky130_fd_sc_hd__nor2_1
X_08288_ input30/X _08341_/B _08342_/A _08344_/A VGND VGND VPWR VPWR _08339_/A sky130_fd_sc_hd__o22a_1
XFILLER_125_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10250_ _10250_/A _10252_/B VGND VGND VPWR VPWR _10250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10181_ _10175_/Y _10179_/Y _10180_/Y VGND VGND VPWR VPWR _10182_/A sky130_fd_sc_hd__o21ai_1
X_13940_ _15392_/A _13940_/B VGND VGND VPWR VPWR _13940_/X sky130_fd_sc_hd__or2_1
XFILLER_59_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15610_ _15539_/Y _15609_/A _15539_/A _15609_/Y _15595_/A VGND VGND VPWR VPWR _16040_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_75_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13871_ _13542_/X _13870_/Y _13542_/X _13870_/Y VGND VGND VPWR VPWR _13873_/B sky130_fd_sc_hd__a2bb2o_1
X_12822_ _12840_/A _12840_/B VGND VGND VPWR VPWR _12822_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15541_ _15536_/Y _15539_/Y _15540_/Y VGND VGND VPWR VPWR _15602_/A sky130_fd_sc_hd__o21ai_2
XFILLER_91_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _12767_/A _12767_/B VGND VGND VPWR VPWR _12753_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11704_ _11677_/X _11703_/X _11677_/X _11703_/X VGND VGND VPWR VPWR _11705_/A sky130_fd_sc_hd__a2bb2oi_4
X_15472_ _12232_/Y _15471_/X _12232_/Y _15471_/X VGND VGND VPWR VPWR _15473_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14423_/A _14423_/B VGND VGND VPWR VPWR _14423_/Y sky130_fd_sc_hd__nor2_1
X_12684_ _12684_/A _12684_/B VGND VGND VPWR VPWR _12684_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11635_ _12863_/A _11636_/B VGND VGND VPWR VPWR _11637_/A sky130_fd_sc_hd__and2_1
XFILLER_11_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14354_ _14380_/A _15950_/A VGND VGND VPWR VPWR _15644_/A sky130_fd_sc_hd__and2_1
X_11566_ _11566_/A _11566_/B VGND VGND VPWR VPWR _11566_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14285_ _12636_/X _14284_/X _12636_/X _14284_/X VGND VGND VPWR VPWR _14285_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13305_ _13305_/A VGND VGND VPWR VPWR _13305_/Y sky130_fd_sc_hd__inv_2
X_10517_ _11833_/A VGND VGND VPWR VPWR _13610_/A sky130_fd_sc_hd__buf_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16024_ _15947_/Y _16023_/X _15947_/Y _16023_/X VGND VGND VPWR VPWR _16030_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13236_ _15066_/A VGND VGND VPWR VPWR _14474_/A sky130_fd_sc_hd__inv_2
X_11497_ _12390_/A VGND VGND VPWR VPWR _12953_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10448_ _11801_/A VGND VGND VPWR VPWR _13519_/A sky130_fd_sc_hd__buf_1
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13167_ _13108_/X _13166_/Y _13108_/X _13166_/Y VGND VGND VPWR VPWR _13190_/B sky130_fd_sc_hd__a2bb2o_1
X_10379_ _11805_/A _10453_/B VGND VGND VPWR VPWR _10379_/Y sky130_fd_sc_hd__nand2_1
X_12118_ _12056_/X _12117_/Y _12056_/X _12117_/Y VGND VGND VPWR VPWR _12145_/B sky130_fd_sc_hd__a2bb2o_1
X_13098_ _14505_/A _13008_/B _13008_/Y VGND VGND VPWR VPWR _13098_/Y sky130_fd_sc_hd__a21oi_1
X_12049_ _12049_/A _12049_/B VGND VGND VPWR VPWR _12049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15808_ _15755_/Y _16197_/A _15807_/Y VGND VGND VPWR VPWR _15808_/X sky130_fd_sc_hd__o21a_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15739_ _14917_/X _15738_/X _14917_/X _15738_/X VGND VGND VPWR VPWR _15740_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_92_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09260_ _10014_/A _08801_/A _10050_/A _09259_/X VGND VGND VPWR VPWR _09260_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09191_ _09429_/A _09191_/B VGND VGND VPWR VPWR _11664_/B sky130_fd_sc_hd__and2_1
XFILLER_119_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08975_ _08901_/X _08973_/X _11378_/B VGND VGND VPWR VPWR _08975_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09527_ _09527_/A _09527_/B VGND VGND VPWR VPWR _09528_/A sky130_fd_sc_hd__or2_1
XFILLER_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09458_ _09458_/A _09458_/B VGND VGND VPWR VPWR _09458_/Y sky130_fd_sc_hd__nor2_1
X_08409_ _08409_/A VGND VGND VPWR VPWR _08409_/Y sky130_fd_sc_hd__inv_2
X_09389_ _09360_/X _09388_/Y _09360_/X _09388_/Y VGND VGND VPWR VPWR _09389_/X sky130_fd_sc_hd__a2bb2o_1
X_11420_ _13405_/A _11420_/B VGND VGND VPWR VPWR _11420_/X sky130_fd_sc_hd__and2_1
XFILLER_61_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11351_ _11351_/A _11350_/X VGND VGND VPWR VPWR _11351_/X sky130_fd_sc_hd__or2b_1
X_10302_ _10455_/A _11225_/A VGND VGND VPWR VPWR _10303_/A sky130_fd_sc_hd__or2_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11282_ _11480_/A VGND VGND VPWR VPWR _14745_/A sky130_fd_sc_hd__buf_1
X_14070_ _11692_/Y _14069_/X _11692_/Y _14069_/X VGND VGND VPWR VPWR _14070_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13021_ _13075_/A _13019_/X _13020_/X VGND VGND VPWR VPWR _13021_/X sky130_fd_sc_hd__o21a_1
X_10233_ _10235_/A _10235_/B VGND VGND VPWR VPWR _10234_/A sky130_fd_sc_hd__or2_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10164_ _10113_/A _10113_/B _10114_/A VGND VGND VPWR VPWR _10167_/A sky130_fd_sc_hd__a21bo_1
XFILLER_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14972_ _14933_/Y _14971_/Y _14961_/Y VGND VGND VPWR VPWR _14972_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10095_ _09954_/Y _10094_/A _09954_/A _10094_/Y VGND VGND VPWR VPWR _11237_/A sky130_fd_sc_hd__a22o_2
X_13923_ _14631_/A _13844_/B _13844_/Y VGND VGND VPWR VPWR _13923_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13854_ _14611_/A _13854_/B VGND VGND VPWR VPWR _13854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12805_ _12775_/A _12775_/B _12775_/Y VGND VGND VPWR VPWR _12805_/Y sky130_fd_sc_hd__o21ai_1
X_15524_ _15524_/A _15524_/B VGND VGND VPWR VPWR _15524_/Y sky130_fd_sc_hd__nand2_1
X_10997_ _11116_/A _10996_/Y _11116_/A _10996_/Y VGND VGND VPWR VPWR _10998_/B sky130_fd_sc_hd__a2bb2o_1
X_13785_ _13541_/X _13784_/Y _13541_/X _13784_/Y VGND VGND VPWR VPWR _13786_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _12690_/A _12690_/B _12690_/Y VGND VGND VPWR VPWR _12736_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15455_ _15455_/A _15455_/B VGND VGND VPWR VPWR _15455_/X sky130_fd_sc_hd__and2_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _10811_/Y _12666_/Y _10683_/Y VGND VGND VPWR VPWR _12668_/A sky130_fd_sc_hd__o21ai_1
X_14406_ _14291_/Y _14404_/X _14405_/Y VGND VGND VPWR VPWR _14406_/X sky130_fd_sc_hd__o21a_1
X_15386_ _15402_/A _15402_/B VGND VGND VPWR VPWR _15462_/A sky130_fd_sc_hd__and2_1
X_11618_ _11620_/A VGND VGND VPWR VPWR _11618_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14337_ _15872_/A _14260_/B _14260_/Y VGND VGND VPWR VPWR _14337_/Y sky130_fd_sc_hd__o21ai_1
X_12598_ _12598_/A VGND VGND VPWR VPWR _12598_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11549_ _12393_/A _11649_/B VGND VGND VPWR VPWR _11549_/Y sky130_fd_sc_hd__nand2_1
X_14268_ _14268_/A VGND VGND VPWR VPWR _14268_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16007_ _16042_/A _16042_/B VGND VGND VPWR VPWR _16007_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14199_ _14112_/A _14112_/B _14112_/Y VGND VGND VPWR VPWR _14199_/X sky130_fd_sc_hd__o21a_1
X_13219_ _13203_/X _13218_/Y _13203_/X _13218_/Y VGND VGND VPWR VPWR _13303_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _10133_/A VGND VGND VPWR VPWR _08760_/Y sky130_fd_sc_hd__inv_2
X_08691_ _08881_/A _08689_/X _08881_/B VGND VGND VPWR VPWR _08691_/X sky130_fd_sc_hd__o21ba_1
XFILLER_81_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09312_ _09313_/A _09313_/B VGND VGND VPWR VPWR _09312_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09243_ _08597_/A _09856_/A _09216_/Y _09242_/X VGND VGND VPWR VPWR _09243_/X sky130_fd_sc_hd__o22a_1
X_09174_ _09757_/A VGND VGND VPWR VPWR _09431_/A sky130_fd_sc_hd__buf_1
XFILLER_119_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08958_ _09538_/A _08635_/A _08637_/A VGND VGND VPWR VPWR _08958_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08889_ _08888_/Y _08864_/X _08888_/Y _08864_/X VGND VGND VPWR VPWR _08978_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10920_ _11018_/A _10917_/X _10919_/X VGND VGND VPWR VPWR _10920_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10851_ _10775_/X _10850_/Y _10775_/X _10850_/Y VGND VGND VPWR VPWR _10919_/B sky130_fd_sc_hd__o2bb2a_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10782_ _10782_/A VGND VGND VPWR VPWR _10782_/Y sky130_fd_sc_hd__inv_2
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _13530_/A _13530_/B _13530_/Y VGND VGND VPWR VPWR _13570_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12521_ _13442_/A _11370_/B _11370_/Y VGND VGND VPWR VPWR _12522_/B sky130_fd_sc_hd__o21a_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A _15240_/B VGND VGND VPWR VPWR _15240_/Y sky130_fd_sc_hd__nand2_1
X_12452_ _12452_/A _12452_/B VGND VGND VPWR VPWR _12452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11403_ _11409_/B _11403_/B VGND VGND VPWR VPWR _12329_/A sky130_fd_sc_hd__or2_1
X_15171_ _15171_/A _15425_/B VGND VGND VPWR VPWR _15171_/Y sky130_fd_sc_hd__nand2_1
X_12383_ _12435_/A _12382_/B _12382_/Y VGND VGND VPWR VPWR _12383_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14122_ _14116_/X _14119_/Y _14876_/A _14121_/Y VGND VGND VPWR VPWR _14122_/X sky130_fd_sc_hd__o22a_1
X_11334_ _11506_/A _11507_/B _11506_/A _11507_/B VGND VGND VPWR VPWR _11334_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14053_ _15461_/A _14032_/B _14032_/X _14052_/X VGND VGND VPWR VPWR _14053_/X sky130_fd_sc_hd__o22a_1
X_11265_ _13371_/A VGND VGND VPWR VPWR _14009_/A sky130_fd_sc_hd__inv_2
XFILLER_79_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13004_ _15146_/A _12920_/B _12920_/Y VGND VGND VPWR VPWR _13004_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10216_ _10216_/A VGND VGND VPWR VPWR _10216_/X sky130_fd_sc_hd__buf_1
XFILLER_121_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11196_ _11090_/X _11195_/X _11090_/X _11195_/X VGND VGND VPWR VPWR _11197_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10147_ _10147_/A _10147_/B VGND VGND VPWR VPWR _10147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14955_ _14952_/Y _14954_/X _14952_/Y _14954_/X VGND VGND VPWR VPWR _14956_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10078_ _10052_/X _10076_/X _10675_/B VGND VGND VPWR VPWR _10078_/X sky130_fd_sc_hd__o21a_1
X_13906_ _13906_/A VGND VGND VPWR VPWR _15410_/A sky130_fd_sc_hd__buf_1
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14886_ _15540_/A _14916_/B VGND VGND VPWR VPWR _14886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13837_ _14644_/A _13838_/B VGND VGND VPWR VPWR _13837_/Y sky130_fd_sc_hd__nor2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13768_ _13813_/A _13766_/X _13767_/X VGND VGND VPWR VPWR _13768_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15507_ _15473_/A _15473_/B _15473_/Y VGND VGND VPWR VPWR _15507_/Y sky130_fd_sc_hd__o21ai_1
X_12719_ _12684_/A _12684_/B _12684_/Y _12718_/X VGND VGND VPWR VPWR _12719_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15438_ _15438_/A _15418_/X VGND VGND VPWR VPWR _15438_/X sky130_fd_sc_hd__or2b_1
X_13699_ _13699_/A _13699_/B VGND VGND VPWR VPWR _13699_/X sky130_fd_sc_hd__or2_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15369_ _15369_/A _15345_/X VGND VGND VPWR VPWR _15369_/X sky130_fd_sc_hd__or2b_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09930_ _09928_/A _09928_/B _09929_/Y VGND VGND VPWR VPWR _09930_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09861_ _09861_/A _09861_/B VGND VGND VPWR VPWR _09924_/A sky130_fd_sc_hd__or2_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08812_ _09217_/A _09455_/B _08715_/X VGND VGND VPWR VPWR _08813_/A sky130_fd_sc_hd__o21ai_1
X_09792_ _09792_/A VGND VGND VPWR VPWR _09793_/B sky130_fd_sc_hd__inv_2
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08743_ _10009_/A _09525_/A VGND VGND VPWR VPWR _08743_/X sky130_fd_sc_hd__or2_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08674_ _09029_/A VGND VGND VPWR VPWR _08674_/Y sky130_fd_sc_hd__inv_2
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09226_ _09801_/A VGND VGND VPWR VPWR _09690_/A sky130_fd_sc_hd__inv_2
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09157_ _08710_/Y _09054_/Y _08740_/X VGND VGND VPWR VPWR _09158_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09088_ _09088_/A VGND VGND VPWR VPWR _09088_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11050_ _12037_/A _10891_/B _10891_/Y VGND VGND VPWR VPWR _11050_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10001_ _09569_/A _09999_/B _09749_/X _10000_/Y VGND VGND VPWR VPWR _10001_/X sky130_fd_sc_hd__o22a_1
XFILLER_1_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14740_ _14780_/A _14738_/X _14739_/X VGND VGND VPWR VPWR _14740_/X sky130_fd_sc_hd__o21a_1
X_11952_ _12994_/A _11895_/B _11895_/Y VGND VGND VPWR VPWR _11952_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14671_ _14597_/A _14597_/B _14594_/X _14597_/Y VGND VGND VPWR VPWR _14671_/X sky130_fd_sc_hd__o2bb2a_1
X_11883_ _11835_/A _11835_/B _11835_/Y VGND VGND VPWR VPWR _11883_/Y sky130_fd_sc_hd__o21ai_1
X_10903_ _10903_/A VGND VGND VPWR VPWR _11411_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16410_ _16406_/Y _16409_/Y _16349_/X _16349_/X _16402_/X VGND VGND VPWR VPWR _16411_/B
+ sky130_fd_sc_hd__o32a_1
X_13622_ _15137_/A _13622_/B VGND VGND VPWR VPWR _13622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10834_ _11007_/A _10951_/B _11007_/A _10951_/B VGND VGND VPWR VPWR _10834_/X sky130_fd_sc_hd__a2bb2o_1
X_16341_ input1/X VGND VGND VPWR VPWR _16361_/A sky130_fd_sc_hd__inv_2
X_13553_ _13553_/A VGND VGND VPWR VPWR _13553_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12504_ _14138_/A VGND VGND VPWR VPWR _13446_/A sky130_fd_sc_hd__buf_1
X_10765_ _11061_/A _11063_/B VGND VGND VPWR VPWR _10765_/X sky130_fd_sc_hd__or2_1
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16272_ _16272_/A VGND VGND VPWR VPWR _16338_/A sky130_fd_sc_hd__buf_1
XFILLER_73_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10696_ _11014_/A _10795_/B _11014_/A _10795_/B VGND VGND VPWR VPWR _10696_/X sky130_fd_sc_hd__a2bb2o_1
X_13484_ _10365_/Y _11750_/A _10316_/Y _13483_/X VGND VGND VPWR VPWR _13484_/X sky130_fd_sc_hd__o22a_1
X_15223_ _15196_/A _15196_/B _15196_/Y _15222_/X VGND VGND VPWR VPWR _15223_/X sky130_fd_sc_hd__a2bb2o_1
X_12435_ _12435_/A _12435_/B VGND VGND VPWR VPWR _12435_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15154_ _15125_/A _15125_/B _15125_/Y _15153_/X VGND VGND VPWR VPWR _15154_/X sky130_fd_sc_hd__a2bb2o_1
X_12366_ _12365_/Y _12258_/X _12281_/Y VGND VGND VPWR VPWR _12366_/X sky130_fd_sc_hd__o21a_1
XFILLER_114_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14105_ _14053_/X _14104_/X _14053_/X _14104_/X VGND VGND VPWR VPWR _14105_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_4_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11317_ _10084_/X _11316_/X _10084_/X _11316_/X VGND VGND VPWR VPWR _11318_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12297_ _14009_/A _12297_/B VGND VGND VPWR VPWR _12297_/Y sky130_fd_sc_hd__nand2_1
X_15085_ _10426_/A _12833_/Y _10422_/A _12830_/X VGND VGND VPWR VPWR _15087_/B sky130_fd_sc_hd__a22o_1
X_14036_ _14036_/A _14036_/B VGND VGND VPWR VPWR _14036_/X sky130_fd_sc_hd__and2_1
X_11248_ _14048_/A _11250_/B VGND VGND VPWR VPWR _11248_/X sky130_fd_sc_hd__and2_1
X_11179_ _14062_/A _11179_/B VGND VGND VPWR VPWR _11179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15987_ _15854_/Y _15986_/X _15854_/Y _15986_/X VGND VGND VPWR VPWR _15987_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_67_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14938_ _15167_/A _14938_/B VGND VGND VPWR VPWR _14938_/Y sky130_fd_sc_hd__nor2_1
X_14869_ _14778_/A _14778_/B _14778_/A _14778_/B VGND VGND VPWR VPWR _14869_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08390_ _08388_/Y _08389_/A _08388_/A _08389_/Y _08303_/A VGND VGND VPWR VPWR _09006_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09011_ _08904_/X _09023_/S _08604_/Y VGND VGND VPWR VPWR _09011_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09913_ _09913_/A _09913_/B VGND VGND VPWR VPWR _10947_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09844_ _09844_/A VGND VGND VPWR VPWR _09844_/Y sky130_fd_sc_hd__inv_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09775_ _09776_/A _09776_/B VGND VGND VPWR VPWR _09775_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08726_ _08717_/A _08717_/B _08717_/X _08725_/Y VGND VGND VPWR VPWR _08726_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08657_ _08657_/A VGND VGND VPWR VPWR _08657_/Y sky130_fd_sc_hd__inv_2
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08588_ _08587_/A _08343_/Y _08587_/Y _08343_/A VGND VGND VPWR VPWR _08589_/B sky130_fd_sc_hd__o22a_1
X_10550_ _10552_/A VGND VGND VPWR VPWR _10550_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10481_ _10436_/X _10480_/X _10436_/X _10480_/X VGND VGND VPWR VPWR _10533_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09209_ _09209_/A _09209_/B VGND VGND VPWR VPWR _09857_/A sky130_fd_sc_hd__or2_2
XFILLER_10_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12220_ _12142_/X _12219_/X _12142_/X _12219_/X VGND VGND VPWR VPWR _12221_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12151_ _13902_/A _12151_/B VGND VGND VPWR VPWR _12151_/X sky130_fd_sc_hd__or2_1
X_11102_ _15057_/A VGND VGND VPWR VPWR _13894_/A sky130_fd_sc_hd__buf_1
X_12082_ _12082_/A _12082_/B VGND VGND VPWR VPWR _12082_/Y sky130_fd_sc_hd__nor2_1
X_15910_ _15910_/A VGND VGND VPWR VPWR _15978_/A sky130_fd_sc_hd__inv_2
XFILLER_110_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11033_ _10913_/X _11032_/X _10913_/X _11032_/X VGND VGND VPWR VPWR _11085_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15841_ _12604_/X _15840_/Y _14232_/B VGND VGND VPWR VPWR _15841_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15772_ _15778_/B _15772_/B VGND VGND VPWR VPWR _16084_/A sky130_fd_sc_hd__or2_1
XFILLER_92_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12984_ _12931_/X _12983_/Y _12931_/X _12983_/Y VGND VGND VPWR VPWR _13020_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14723_ _13937_/X _14721_/Y _14722_/Y VGND VGND VPWR VPWR _14723_/X sky130_fd_sc_hd__o21a_1
X_11935_ _11910_/X _11934_/Y _11910_/X _11934_/Y VGND VGND VPWR VPWR _11978_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14654_ _15339_/A _14654_/B VGND VGND VPWR VPWR _14654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13605_ _13575_/Y _13604_/Y _13575_/Y _13604_/Y VGND VGND VPWR VPWR _13606_/B sky130_fd_sc_hd__a2bb2o_1
X_11866_ _11846_/X _11865_/X _11846_/X _11865_/X VGND VGND VPWR VPWR _11909_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14585_ _14547_/Y _14583_/X _14584_/Y VGND VGND VPWR VPWR _14585_/X sky130_fd_sc_hd__o21a_1
X_11797_ _13560_/A _11770_/B _11770_/X _11796_/X VGND VGND VPWR VPWR _11797_/X sky130_fd_sc_hd__o22a_1
X_10817_ _10242_/B _10155_/B _10155_/Y VGND VGND VPWR VPWR _10818_/A sky130_fd_sc_hd__a21oi_1
X_16324_ _16324_/A _16324_/B VGND VGND VPWR VPWR _16324_/Y sky130_fd_sc_hd__nand2_1
X_13536_ _15036_/A _13519_/B _13519_/Y _13535_/X VGND VGND VPWR VPWR _13536_/X sky130_fd_sc_hd__a2bb2o_1
X_10748_ _09952_/A _09631_/B _09632_/A VGND VGND VPWR VPWR _10749_/A sky130_fd_sc_hd__o21ai_1
X_16255_ _16255_/A _16255_/B VGND VGND VPWR VPWR _16255_/Y sky130_fd_sc_hd__nand2_1
X_13467_ _12425_/A _12679_/B _12679_/Y _12720_/X VGND VGND VPWR VPWR _13467_/Y sky130_fd_sc_hd__o2bb2ai_1
X_15206_ _15140_/A _15140_/B _15140_/Y VGND VGND VPWR VPWR _15206_/Y sky130_fd_sc_hd__o21ai_1
X_12418_ _12682_/A _12417_/B _12417_/X _12379_/B VGND VGND VPWR VPWR _12419_/B sky130_fd_sc_hd__a22o_1
X_10679_ _10243_/B _10159_/B _10159_/Y VGND VGND VPWR VPWR _10680_/A sky130_fd_sc_hd__a21oi_1
X_16186_ _16262_/A _16328_/A VGND VGND VPWR VPWR _16186_/Y sky130_fd_sc_hd__nor2_1
X_13398_ _15524_/A VGND VGND VPWR VPWR _14093_/A sky130_fd_sc_hd__inv_2
XFILLER_126_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12349_ _12349_/A _12349_/B VGND VGND VPWR VPWR _12349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15137_ _15137_/A _15137_/B VGND VGND VPWR VPWR _15137_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15068_ _15037_/X _15067_/X _15037_/X _15067_/X VGND VGND VPWR VPWR _15069_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14019_ _15410_/A _13952_/B _13952_/Y VGND VGND VPWR VPWR _14019_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09560_ _08694_/A _09152_/A _09526_/Y _09559_/X VGND VGND VPWR VPWR _09560_/X sky130_fd_sc_hd__o22a_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09491_ _08798_/X _09468_/X _08798_/X _09468_/X VGND VGND VPWR VPWR _09492_/B sky130_fd_sc_hd__o2bb2a_1
X_08511_ _08567_/B VGND VGND VPWR VPWR _09791_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08442_ _08440_/A _08323_/Y _08440_/Y _08323_/A _08441_/X VGND VGND VPWR VPWR _08554_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08373_ input17/X _08254_/B _08327_/B _08434_/A VGND VGND VPWR VPWR _08440_/A sky130_fd_sc_hd__o22a_1
XFILLER_129_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ _09808_/A _09503_/B _09817_/A _09817_/B _09826_/X VGND VGND VPWR VPWR _09827_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09758_ _09739_/A _09739_/B _09742_/A VGND VGND VPWR VPWR _10043_/A sky130_fd_sc_hd__a21bo_1
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08709_ _09331_/A _09476_/B VGND VGND VPWR VPWR _08709_/Y sky130_fd_sc_hd__nor2_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11720_/A _11720_/B VGND VGND VPWR VPWR _11731_/B sky130_fd_sc_hd__or2_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09689_ _09689_/A _09689_/B VGND VGND VPWR VPWR _09692_/A sky130_fd_sc_hd__or2_1
XFILLER_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11648_/X _11650_/X _11648_/X _11650_/X VGND VGND VPWR VPWR _11654_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14370_ _14370_/A VGND VGND VPWR VPWR _15662_/B sky130_fd_sc_hd__inv_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10602_ _10602_/A VGND VGND VPWR VPWR _10602_/Y sky130_fd_sc_hd__inv_2
X_11582_ _09440_/X _11581_/X _09440_/X _11581_/X VGND VGND VPWR VPWR _11583_/B sky130_fd_sc_hd__a2bb2o_1
X_13321_ _13296_/A _13320_/Y _13296_/A _13320_/Y VGND VGND VPWR VPWR _13367_/B sky130_fd_sc_hd__a2bb2o_1
X_10533_ _11843_/A _10533_/B VGND VGND VPWR VPWR _10533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _16040_/A _16040_/B VGND VGND VPWR VPWR _16040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13252_ _14423_/A VGND VGND VPWR VPWR _14729_/A sky130_fd_sc_hd__buf_1
XFILLER_10_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10464_ _10462_/A _10461_/Y _10462_/Y _10461_/A _10974_/A VGND VGND VPWR VPWR _10554_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_123_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12203_ _14012_/A _12203_/B VGND VGND VPWR VPWR _12203_/Y sky130_fd_sc_hd__nand2_1
X_13183_ _15329_/A _13182_/B _12043_/Y _13182_/Y VGND VGND VPWR VPWR _13183_/X sky130_fd_sc_hd__o2bb2a_1
X_10395_ _09286_/Y _10394_/A _09286_/A _10394_/Y _09392_/A VGND VGND VPWR VPWR _10396_/A
+ sky130_fd_sc_hd__o221a_1
X_12134_ _12135_/A _12135_/B VGND VGND VPWR VPWR _12134_/X sky130_fd_sc_hd__or2_1
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12065_ _12104_/A VGND VGND VPWR VPWR _13200_/A sky130_fd_sc_hd__buf_1
XFILLER_77_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11016_ _12850_/A VGND VGND VPWR VPWR _15066_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15824_ _15706_/X _15822_/X _15834_/B VGND VGND VPWR VPWR _15824_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15755_ _16106_/A _15807_/B VGND VGND VPWR VPWR _15755_/Y sky130_fd_sc_hd__nor2_1
X_12967_ _14600_/A _12940_/B _12940_/Y VGND VGND VPWR VPWR _12967_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15686_ _15585_/Y _15684_/X _15685_/Y VGND VGND VPWR VPWR _15694_/A sky130_fd_sc_hd__o21a_1
X_14706_ _15337_/A _14652_/B _14652_/Y VGND VGND VPWR VPWR _14706_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12898_ _12843_/X _12897_/Y _12843_/X _12897_/Y VGND VGND VPWR VPWR _12930_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11918_ _11918_/A _11918_/B VGND VGND VPWR VPWR _11918_/X sky130_fd_sc_hd__or2_1
X_14637_ _14575_/X _14636_/Y _14575_/X _14636_/Y VGND VGND VPWR VPWR _14648_/B sky130_fd_sc_hd__a2bb2o_1
X_11849_ _11847_/A _11847_/B _11847_/X _11848_/Y VGND VGND VPWR VPWR _11913_/B sky130_fd_sc_hd__a22o_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _14568_/A VGND VGND VPWR VPWR _15270_/A sky130_fd_sc_hd__buf_1
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16307_ _16252_/X _16306_/Y _16252_/X _16306_/Y VGND VGND VPWR VPWR _16320_/B sky130_fd_sc_hd__o2bb2a_1
X_14499_ _14460_/X _14498_/Y _14460_/X _14498_/Y VGND VGND VPWR VPWR _14512_/B sky130_fd_sc_hd__a2bb2o_1
X_13519_ _13519_/A _13519_/B VGND VGND VPWR VPWR _13519_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16238_ _16238_/A _16238_/B VGND VGND VPWR VPWR _16249_/B sky130_fd_sc_hd__or2_1
X_16169_ _16266_/B VGND VGND VPWR VPWR _16332_/A sky130_fd_sc_hd__buf_1
XFILLER_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08991_ _09478_/A VGND VGND VPWR VPWR _09518_/A sky130_fd_sc_hd__buf_1
XFILLER_96_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09612_ _09977_/A VGND VGND VPWR VPWR _09978_/A sky130_fd_sc_hd__buf_1
XFILLER_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09543_ _09540_/A _09540_/B _09540_/X _09628_/B VGND VGND VPWR VPWR _09543_/X sky130_fd_sc_hd__a22o_1
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09474_ _10010_/A _09474_/B VGND VGND VPWR VPWR _09474_/X sky130_fd_sc_hd__or2_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08425_ _08424_/A _08338_/Y _08424_/Y _08338_/A _08441_/A VGND VGND VPWR VPWR _09213_/A
+ sky130_fd_sc_hd__o221a_1
X_08356_ _08354_/Y _08355_/A _08354_/A _08355_/Y _08303_/A VGND VGND VPWR VPWR _09225_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08287_ input29/X _08346_/B _08347_/A _08349_/A VGND VGND VPWR VPWR _08344_/A sky130_fd_sc_hd__o22a_1
XFILLER_124_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10180_ _10180_/A _10180_/B VGND VGND VPWR VPWR _10180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13870_ _15104_/A _13498_/B _13498_/Y VGND VGND VPWR VPWR _13870_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12821_ _12764_/X _12820_/Y _12764_/X _12820_/Y VGND VGND VPWR VPWR _12840_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15540_ _15540_/A _15540_/B VGND VGND VPWR VPWR _15540_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12752_ _12710_/X _12751_/X _12710_/X _12751_/X VGND VGND VPWR VPWR _12767_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15471_ _15471_/A _15395_/X VGND VGND VPWR VPWR _15471_/X sky130_fd_sc_hd__or2b_1
X_11703_ _11688_/Y _11702_/Y _11688_/Y _11702_/Y VGND VGND VPWR VPWR _11703_/X sky130_fd_sc_hd__a2bb2o_2
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _11326_/A _12674_/A _11326_/Y _12674_/Y VGND VGND VPWR VPWR _12684_/B sky130_fd_sc_hd__o22a_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14422_ _11768_/Y _14418_/X _11768_/Y _14418_/X VGND VGND VPWR VPWR _14423_/B sky130_fd_sc_hd__o2bb2a_1
X_11634_ _11630_/X _11633_/X _11630_/X _11633_/X VGND VGND VPWR VPWR _11636_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14353_ _14353_/A _14353_/B VGND VGND VPWR VPWR _15950_/A sky130_fd_sc_hd__or2_1
X_11565_ _13448_/A _11564_/B _11564_/Y VGND VGND VPWR VPWR _11566_/B sky130_fd_sc_hd__o21a_1
XFILLER_11_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14284_ _14284_/A _12637_/X VGND VGND VPWR VPWR _14284_/X sky130_fd_sc_hd__or2b_1
X_13304_ _13220_/Y _13302_/Y _13303_/Y VGND VGND VPWR VPWR _13305_/A sky130_fd_sc_hd__o21ai_1
X_11496_ _11590_/A _11496_/B VGND VGND VPWR VPWR _12390_/A sky130_fd_sc_hd__or2_1
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10516_ _09403_/X _08931_/Y _08931_/A _10515_/Y _11592_/A VGND VGND VPWR VPWR _11833_/A
+ sky130_fd_sc_hd__a221o_2
X_16023_ _16023_/A _15948_/X VGND VGND VPWR VPWR _16023_/X sky130_fd_sc_hd__or2b_1
XFILLER_108_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13235_ _14737_/A _13294_/B VGND VGND VPWR VPWR _13235_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10447_ _09970_/A _10445_/Y _09970_/Y _10445_/A _10957_/A VGND VGND VPWR VPWR _11801_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13166_ _15258_/A _13109_/B _13109_/Y VGND VGND VPWR VPWR _13166_/Y sky130_fd_sc_hd__o21ai_1
X_10378_ _10377_/A _10376_/Y _10377_/Y _10376_/A _10463_/A VGND VGND VPWR VPWR _10453_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13097_ _13101_/A VGND VGND VPWR VPWR _14568_/A sky130_fd_sc_hd__buf_1
X_12117_ _13192_/A _12057_/B _12057_/Y VGND VGND VPWR VPWR _12117_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12048_ _12043_/Y _12046_/Y _12047_/Y VGND VGND VPWR VPWR _12048_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15807_ _16106_/A _15807_/B VGND VGND VPWR VPWR _15807_/Y sky130_fd_sc_hd__nand2_1
X_13999_ _15425_/A _13972_/A _13973_/Y _13998_/Y VGND VGND VPWR VPWR _13999_/X sky130_fd_sc_hd__o22a_1
X_15738_ _15542_/A _14918_/B _14918_/Y VGND VGND VPWR VPWR _15738_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15669_ _15669_/A _15669_/B VGND VGND VPWR VPWR _15669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09190_ _11664_/A _09190_/B VGND VGND VPWR VPWR _09190_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08974_ _08974_/A _08974_/B VGND VGND VPWR VPWR _11378_/B sky130_fd_sc_hd__or2_1
XFILLER_130_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09526_ _09526_/A VGND VGND VPWR VPWR _09526_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09457_ _09498_/A _09457_/B VGND VGND VPWR VPWR _09457_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08408_ _09228_/A _08386_/Y _08407_/Y VGND VGND VPWR VPWR _08408_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_51_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09388_ _09429_/B _11574_/A _09365_/X _11576_/A VGND VGND VPWR VPWR _09388_/Y sky130_fd_sc_hd__a22oi_1
X_08339_ _08339_/A VGND VGND VPWR VPWR _08339_/Y sky130_fd_sc_hd__inv_2
X_11350_ _13890_/A _11350_/B VGND VGND VPWR VPWR _11350_/X sky130_fd_sc_hd__or2_1
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10301_ _09112_/A _10300_/X _09112_/A _10300_/X VGND VGND VPWR VPWR _11225_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_118_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11281_ _12290_/A VGND VGND VPWR VPWR _11480_/A sky130_fd_sc_hd__inv_2
X_13020_ _14485_/A _13020_/B VGND VGND VPWR VPWR _13020_/X sky130_fd_sc_hd__or2_1
XFILLER_121_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10232_ _09298_/A _10230_/B _10231_/Y _10108_/Y VGND VGND VPWR VPWR _10235_/B sky130_fd_sc_hd__o22a_1
XFILLER_121_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10163_ _10163_/A _10163_/B VGND VGND VPWR VPWR _10163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14971_ _14971_/A _14971_/B VGND VGND VPWR VPWR _14971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10094_ _10094_/A VGND VGND VPWR VPWR _10094_/Y sky130_fd_sc_hd__inv_2
X_13922_ _13922_/A VGND VGND VPWR VPWR _15402_/A sky130_fd_sc_hd__buf_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13853_ _13812_/Y _13851_/X _13852_/Y VGND VGND VPWR VPWR _13853_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12804_ _12852_/A _12852_/B VGND VGND VPWR VPWR _12804_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15523_ _15476_/X _15522_/Y _15476_/X _15522_/Y VGND VGND VPWR VPWR _15632_/A sky130_fd_sc_hd__a2bb2o_1
X_10996_ _13703_/A _11115_/B _10995_/Y VGND VGND VPWR VPWR _10996_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13784_ _15051_/A _13501_/B _13501_/Y VGND VGND VPWR VPWR _13784_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12779_/A _12779_/B VGND VGND VPWR VPWR _12735_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15454_ _15407_/X _15453_/X _15407_/X _15453_/X VGND VGND VPWR VPWR _15455_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12666_ _12666_/A VGND VGND VPWR VPWR _12666_/Y sky130_fd_sc_hd__inv_2
X_14405_ _15982_/A _14405_/B VGND VGND VPWR VPWR _14405_/Y sky130_fd_sc_hd__nand2_1
X_12597_ _14906_/A _11422_/B _11422_/Y VGND VGND VPWR VPWR _12598_/A sky130_fd_sc_hd__a21oi_1
X_15385_ _15334_/X _15384_/X _15334_/X _15384_/X VGND VGND VPWR VPWR _15402_/B sky130_fd_sc_hd__a2bb2o_1
X_11617_ _12679_/A _11616_/B _11616_/Y VGND VGND VPWR VPWR _11617_/Y sky130_fd_sc_hd__a21oi_1
X_14336_ _14386_/A _15956_/A VGND VGND VPWR VPWR _15620_/A sky130_fd_sc_hd__and2_1
X_11548_ _11493_/X _11547_/Y _11493_/X _11547_/Y VGND VGND VPWR VPWR _11649_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14267_ _14204_/Y _14265_/Y _14266_/Y VGND VGND VPWR VPWR _14268_/A sky130_fd_sc_hd__o21ai_1
X_11479_ _15107_/A VGND VGND VPWR VPWR _13545_/A sky130_fd_sc_hd__buf_1
X_16006_ _15959_/X _16005_/X _15959_/X _16005_/X VGND VGND VPWR VPWR _16042_/B sky130_fd_sc_hd__a2bb2o_1
X_14198_ _15863_/A _14269_/B VGND VGND VPWR VPWR _14198_/Y sky130_fd_sc_hd__nor2_1
X_13218_ _13204_/A _13204_/B _13204_/Y VGND VGND VPWR VPWR _13218_/Y sky130_fd_sc_hd__o21ai_1
X_13149_ _13120_/X _13148_/Y _13120_/X _13148_/Y VGND VGND VPWR VPWR _13202_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08690_ _08690_/A _10118_/B VGND VGND VPWR VPWR _08881_/B sky130_fd_sc_hd__and2_1
XFILLER_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09311_ _09946_/A _09309_/Y _09310_/Y VGND VGND VPWR VPWR _09313_/B sky130_fd_sc_hd__o21ai_1
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09242_ _08610_/A _09803_/A _09220_/Y _09241_/X VGND VGND VPWR VPWR _09242_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09173_ _10010_/B _09165_/B _09166_/B VGND VGND VPWR VPWR _09757_/A sky130_fd_sc_hd__a21bo_1
XFILLER_130_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08957_ _08960_/A _08960_/B VGND VGND VPWR VPWR _08957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08888_ _09470_/A _08786_/B _08786_/Y VGND VGND VPWR VPWR _08888_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10850_ _13063_/A _10704_/B _10704_/Y VGND VGND VPWR VPWR _10850_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10781_ _11978_/A _10781_/B VGND VGND VPWR VPWR _10781_/Y sky130_fd_sc_hd__nor2_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09509_ _09498_/A _09498_/B _09498_/Y _09508_/X VGND VGND VPWR VPWR _09509_/X sky130_fd_sc_hd__o2bb2a_1
X_12520_ _14126_/A VGND VGND VPWR VPWR _13442_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12448_/X _12450_/X _12448_/X _12450_/X VGND VGND VPWR VPWR _12452_/B sky130_fd_sc_hd__a2bb2o_1
X_15170_ _15168_/X _15169_/Y _15168_/X _15169_/Y VGND VGND VPWR VPWR _15425_/B sky130_fd_sc_hd__a2bb2o_1
X_11402_ _08951_/Y _11401_/X _08951_/Y _11401_/X VGND VGND VPWR VPWR _11403_/B sky130_fd_sc_hd__a2bb2oi_2
X_14121_ _14121_/A VGND VGND VPWR VPWR _14121_/Y sky130_fd_sc_hd__inv_2
X_12382_ _12435_/A _12382_/B VGND VGND VPWR VPWR _12382_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11333_ _11313_/X _11332_/X _11313_/X _11332_/X VGND VGND VPWR VPWR _11507_/B sky130_fd_sc_hd__a2bb2o_1
X_14052_ _15464_/A _14036_/B _14036_/X _14051_/X VGND VGND VPWR VPWR _14052_/X sky130_fd_sc_hd__o22a_1
X_11264_ _09179_/Y _11263_/A _09179_/A _11263_/Y _09204_/X VGND VGND VPWR VPWR _13371_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13003_ _13003_/A VGND VGND VPWR VPWR _15146_/A sky130_fd_sc_hd__buf_1
X_10215_ _10215_/A VGND VGND VPWR VPWR _10455_/A sky130_fd_sc_hd__clkbuf_2
X_11195_ _11195_/A _11091_/X VGND VGND VPWR VPWR _11195_/X sky130_fd_sc_hd__or2b_1
XFILLER_79_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10146_ _08778_/B _10131_/B _10132_/B VGND VGND VPWR VPWR _10147_/B sky130_fd_sc_hd__a21bo_1
X_14954_ _14834_/X _14953_/Y _14851_/Y VGND VGND VPWR VPWR _14954_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10077_ _10077_/A _10077_/B VGND VGND VPWR VPWR _10675_/B sky130_fd_sc_hd__or2_1
X_13905_ _15412_/A _13954_/B VGND VGND VPWR VPWR _13905_/Y sky130_fd_sc_hd__nor2_1
X_14885_ _14821_/X _14884_/X _14821_/X _14884_/X VGND VGND VPWR VPWR _14916_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13836_ _13755_/A _13835_/Y _13755_/A _13835_/Y VGND VGND VPWR VPWR _13838_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13767_ _13767_/A _13767_/B VGND VGND VPWR VPWR _13767_/X sky130_fd_sc_hd__or2_1
XFILLER_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10979_ _10965_/X _10978_/Y _10965_/X _10978_/Y VGND VGND VPWR VPWR _11138_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_16_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15506_ _15542_/A _15542_/B VGND VGND VPWR VPWR _15600_/A sky130_fd_sc_hd__and2_1
X_12718_ _12686_/A _12686_/B _12686_/Y _12717_/X VGND VGND VPWR VPWR _12718_/X sky130_fd_sc_hd__o2bb2a_1
X_15437_ _15437_/A _15437_/B VGND VGND VPWR VPWR _15437_/X sky130_fd_sc_hd__and2_1
X_13698_ _13733_/A _13696_/X _13697_/X VGND VGND VPWR VPWR _13698_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12649_ _12650_/A _12650_/B VGND VGND VPWR VPWR _12649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15368_ _15414_/A _15414_/B VGND VGND VPWR VPWR _15444_/A sky130_fd_sc_hd__and2_1
XFILLER_116_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14319_ _13438_/A _13438_/B _13438_/Y VGND VGND VPWR VPWR _14319_/X sky130_fd_sc_hd__o21a_1
X_15299_ _15349_/A _15349_/B VGND VGND VPWR VPWR _15363_/A sky130_fd_sc_hd__and2_1
XFILLER_116_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09860_ _09860_/A _09914_/A VGND VGND VPWR VPWR _09861_/B sky130_fd_sc_hd__or2_1
XFILLER_124_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08811_ _09456_/A VGND VGND VPWR VPWR _09496_/A sky130_fd_sc_hd__buf_1
X_09791_ _09791_/A _09791_/B _09791_/C VGND VGND VPWR VPWR _09792_/A sky130_fd_sc_hd__or3_2
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08742_ _08742_/A VGND VGND VPWR VPWR _08742_/Y sky130_fd_sc_hd__inv_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08673_ _10228_/A _10098_/A VGND VGND VPWR VPWR _09029_/A sky130_fd_sc_hd__or2_1
XFILLER_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09225_ _09225_/A _09225_/B VGND VGND VPWR VPWR _09801_/A sky130_fd_sc_hd__or2_1
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09156_ _09525_/B _09156_/B VGND VGND VPWR VPWR _09156_/X sky130_fd_sc_hd__or2_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09087_ _09551_/B _09034_/B _09035_/B VGND VGND VPWR VPWR _09088_/A sky130_fd_sc_hd__a21bo_1
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10000_ _10000_/A VGND VGND VPWR VPWR _10000_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09989_ _09989_/A _09990_/B VGND VGND VPWR VPWR _09989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11951_ _13083_/A _11968_/B VGND VGND VPWR VPWR _11951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10902_ _10765_/X _10901_/X _10765_/X _10901_/X VGND VGND VPWR VPWR _10907_/B sky130_fd_sc_hd__a2bb2o_1
X_11882_ _12994_/A _11895_/B VGND VGND VPWR VPWR _11882_/Y sky130_fd_sc_hd__nor2_1
X_14670_ _14600_/A _14600_/B _14593_/X _14600_/Y VGND VGND VPWR VPWR _14670_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13621_ _13621_/A VGND VGND VPWR VPWR _15137_/A sky130_fd_sc_hd__buf_1
X_10833_ _10802_/X _10832_/X _10802_/X _10832_/X VGND VGND VPWR VPWR _10951_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16340_ _16278_/X _16339_/X _16278_/X _16339_/X VGND VGND VPWR VPWR _16392_/A sky130_fd_sc_hd__a2bb2o_1
X_10764_ _10764_/A _13006_/A VGND VGND VPWR VPWR _11063_/B sky130_fd_sc_hd__nand2_1
X_13552_ _13552_/A _13552_/B VGND VGND VPWR VPWR _13553_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12503_ _12639_/A _12639_/B VGND VGND VPWR VPWR _14171_/A sky130_fd_sc_hd__and2_1
XFILLER_40_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16271_ _16154_/Y _16269_/X _16270_/Y VGND VGND VPWR VPWR _16271_/X sky130_fd_sc_hd__o21a_1
X_10695_ _10664_/X _10694_/X _10664_/X _10694_/X VGND VGND VPWR VPWR _10795_/B sky130_fd_sc_hd__a2bb2o_1
X_13483_ _10296_/A _12701_/A _10325_/Y _13482_/X VGND VGND VPWR VPWR _13483_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15222_ _15199_/A _15199_/B _15199_/Y _15221_/X VGND VGND VPWR VPWR _15222_/X sky130_fd_sc_hd__a2bb2o_1
X_12434_ _12435_/A VGND VGND VPWR VPWR _12785_/A sky130_fd_sc_hd__buf_1
X_15153_ _15128_/A _15128_/B _15128_/Y _15152_/X VGND VGND VPWR VPWR _15153_/X sky130_fd_sc_hd__a2bb2o_1
X_12365_ _12365_/A _12365_/B VGND VGND VPWR VPWR _12365_/Y sky130_fd_sc_hd__nor2_1
X_14104_ _15458_/A _14028_/B _14028_/A _14028_/B VGND VGND VPWR VPWR _14104_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15084_ _15084_/A _15084_/B VGND VGND VPWR VPWR _15084_/Y sky130_fd_sc_hd__nand2_1
X_11316_ _10040_/X _11316_/B VGND VGND VPWR VPWR _11316_/X sky130_fd_sc_hd__and2b_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14035_ _13943_/X _14034_/Y _13943_/X _14034_/Y VGND VGND VPWR VPWR _14036_/B sky130_fd_sc_hd__a2bb2o_1
X_12296_ _12248_/X _12295_/X _12248_/X _12295_/X VGND VGND VPWR VPWR _12297_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11247_ _11245_/X _11246_/X _11245_/X _11246_/X VGND VGND VPWR VPWR _11250_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11178_ _11094_/X _11177_/X _11094_/X _11177_/X VGND VGND VPWR VPWR _11179_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10129_ _10129_/A _10129_/B VGND VGND VPWR VPWR _10130_/B sky130_fd_sc_hd__or2_1
X_15986_ _15983_/Y _15985_/X _15983_/Y _15985_/X VGND VGND VPWR VPWR _15986_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14937_ _12437_/A _14936_/X _12437_/A _14936_/X VGND VGND VPWR VPWR _14938_/B sky130_fd_sc_hd__o2bb2a_1
X_14868_ _14868_/A VGND VGND VPWR VPWR _15548_/A sky130_fd_sc_hd__buf_1
XFILLER_63_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13819_ _13819_/A _13763_/X VGND VGND VPWR VPWR _13819_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14799_ _15461_/A VGND VGND VPWR VPWR _14802_/A sky130_fd_sc_hd__buf_1
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16469_ _08229_/A _16469_/D VGND VGND VPWR VPWR _16469_/Q sky130_fd_sc_hd__dfxtp_1
X_09010_ _09496_/A _09024_/S _09221_/B VGND VGND VPWR VPWR _09023_/S sky130_fd_sc_hd__a21oi_1
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09912_ _09913_/A _09913_/B VGND VGND VPWR VPWR _10947_/B sky130_fd_sc_hd__and2_1
XFILLER_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09843_ _09843_/A _09843_/B VGND VGND VPWR VPWR _10491_/B sky130_fd_sc_hd__nor2_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09774_ _10077_/A _09772_/Y _09773_/Y VGND VGND VPWR VPWR _09776_/B sky130_fd_sc_hd__o21ai_1
X_08725_ _08718_/Y _08723_/X _08724_/X VGND VGND VPWR VPWR _08725_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08656_ _08656_/A _09684_/A VGND VGND VPWR VPWR _08657_/A sky130_fd_sc_hd__or2_1
XFILLER_27_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08587_ _08587_/A VGND VGND VPWR VPWR _08587_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09208_ _14062_/A VGND VGND VPWR VPWR _15443_/A sky130_fd_sc_hd__buf_1
X_10480_ _10441_/X _10538_/B _10441_/X _10538_/B VGND VGND VPWR VPWR _10480_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09139_ _09531_/B _09037_/B _09038_/B VGND VGND VPWR VPWR _09140_/A sky130_fd_sc_hd__a21bo_1
XFILLER_118_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12150_ _12210_/A _12148_/X _12149_/X VGND VGND VPWR VPWR _12150_/X sky130_fd_sc_hd__o21a_1
X_11101_ _12856_/A VGND VGND VPWR VPWR _15057_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12081_ _12080_/A _12080_/B _12080_/X _11997_/B VGND VGND VPWR VPWR _12172_/B sky130_fd_sc_hd__a22o_1
XFILLER_1_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11032_ _10867_/A _10867_/B _10867_/A _10867_/B VGND VGND VPWR VPWR _11032_/X sky130_fd_sc_hd__a2bb2o_1
X_15840_ _15840_/A VGND VGND VPWR VPWR _15840_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15771_ _12610_/A _15770_/A _12610_/Y _15770_/Y VGND VGND VPWR VPWR _15772_/B sky130_fd_sc_hd__o22a_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12983_ _14467_/A _12932_/B _12932_/Y VGND VGND VPWR VPWR _12983_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14722_ _14722_/A _14722_/B VGND VGND VPWR VPWR _14722_/Y sky130_fd_sc_hd__nand2_1
X_11934_ _13637_/A _11981_/B _11933_/Y VGND VGND VPWR VPWR _11934_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14653_ _14630_/Y _14651_/X _14652_/Y VGND VGND VPWR VPWR _14653_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13604_ _13568_/A _13568_/B _13569_/A VGND VGND VPWR VPWR _13604_/Y sky130_fd_sc_hd__o21ai_1
X_11865_ _10543_/X _11911_/B _10543_/X _11911_/B VGND VGND VPWR VPWR _11865_/X sky130_fd_sc_hd__a2bb2o_1
X_14584_ _14584_/A _14584_/B VGND VGND VPWR VPWR _14584_/Y sky130_fd_sc_hd__nand2_1
X_11796_ _13564_/A _11775_/B _11775_/X _11795_/X VGND VGND VPWR VPWR _11796_/X sky130_fd_sc_hd__o22a_1
X_10816_ _10816_/A VGND VGND VPWR VPWR _12082_/A sky130_fd_sc_hd__inv_2
XFILLER_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16323_ _16305_/Y _16321_/X _16322_/Y VGND VGND VPWR VPWR _16323_/X sky130_fd_sc_hd__o21a_1
X_10747_ _13088_/A _10747_/B VGND VGND VPWR VPWR _10747_/Y sky130_fd_sc_hd__nand2_1
X_13535_ _15034_/A _13522_/B _13522_/Y _13534_/X VGND VGND VPWR VPWR _13535_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16254_ _16221_/Y _16252_/X _16253_/Y VGND VGND VPWR VPWR _16254_/X sky130_fd_sc_hd__o21a_1
X_13466_ _13461_/Y _13465_/Y _13461_/Y _13465_/Y VGND VGND VPWR VPWR _13466_/X sky130_fd_sc_hd__a2bb2o_1
X_10678_ _10678_/A VGND VGND VPWR VPWR _11992_/A sky130_fd_sc_hd__inv_2
XFILLER_126_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15205_ _15205_/A _15205_/B VGND VGND VPWR VPWR _15205_/Y sky130_fd_sc_hd__nand2_1
X_12417_ _12682_/A _12417_/B VGND VGND VPWR VPWR _12417_/X sky130_fd_sc_hd__or2_1
X_16185_ _16262_/B VGND VGND VPWR VPWR _16328_/A sky130_fd_sc_hd__buf_1
X_13397_ _14098_/A VGND VGND VPWR VPWR _14101_/A sky130_fd_sc_hd__buf_1
XFILLER_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12348_ _12242_/X _12347_/Y _12242_/X _12347_/Y VGND VGND VPWR VPWR _12549_/A sky130_fd_sc_hd__a2bb2o_1
X_15136_ _15090_/X _15135_/Y _15090_/X _15135_/Y VGND VGND VPWR VPWR _15137_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15067_ _15067_/A _15038_/X VGND VGND VPWR VPWR _15067_/X sky130_fd_sc_hd__or2b_1
X_12279_ _11273_/A _12367_/B _11273_/A _12367_/B VGND VGND VPWR VPWR _12279_/X sky130_fd_sc_hd__a2bb2o_1
X_14018_ _14018_/A _14058_/B VGND VGND VPWR VPWR _14117_/A sky130_fd_sc_hd__and2_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15969_ _15966_/A _15966_/B _15966_/Y _15968_/X VGND VGND VPWR VPWR _15969_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_82_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09490_ _09490_/A _09490_/B VGND VGND VPWR VPWR _09490_/Y sky130_fd_sc_hd__nor2_1
X_08510_ _08656_/A VGND VGND VPWR VPWR _08567_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08441_ _08441_/A VGND VGND VPWR VPWR _08441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08372_ input16/X _08257_/B _08332_/B _08429_/A VGND VGND VPWR VPWR _08434_/A sky130_fd_sc_hd__o22a_1
XFILLER_117_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ _09826_/A _09826_/B VGND VGND VPWR VPWR _09826_/X sky130_fd_sc_hd__or2_1
XFILLER_104_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09757_ _09757_/A VGND VGND VPWR VPWR _09785_/A sky130_fd_sc_hd__inv_2
X_08708_ _09448_/A _08755_/A VGND VGND VPWR VPWR _08708_/Y sky130_fd_sc_hd__nor2_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09688_ _08632_/X _09690_/B _08632_/X _09690_/B VGND VGND VPWR VPWR _09689_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08639_ _08660_/A _08639_/B VGND VGND VPWR VPWR _09459_/B sky130_fd_sc_hd__or2_2
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11649_/Y _11486_/Y _11549_/Y VGND VGND VPWR VPWR _11650_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11581_ _09169_/A _09363_/A _09429_/X VGND VGND VPWR VPWR _11581_/X sky130_fd_sc_hd__o21a_1
X_10601_ _09714_/A _09714_/B _09714_/Y VGND VGND VPWR VPWR _10602_/A sky130_fd_sc_hd__a21oi_1
X_13320_ _14739_/A _13297_/B _13297_/Y VGND VGND VPWR VPWR _13320_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10532_ _10489_/Y _10530_/X _10531_/Y VGND VGND VPWR VPWR _10532_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13251_ _15075_/A VGND VGND VPWR VPWR _14423_/A sky130_fd_sc_hd__inv_2
X_10463_ _10463_/A VGND VGND VPWR VPWR _10974_/A sky130_fd_sc_hd__clkbuf_2
X_13182_ _13833_/A _13182_/B VGND VGND VPWR VPWR _13182_/Y sky130_fd_sc_hd__nor2_1
X_12202_ _12154_/X _12201_/X _12154_/X _12201_/X VGND VGND VPWR VPWR _12203_/B sky130_fd_sc_hd__a2bb2o_1
X_10394_ _10394_/A VGND VGND VPWR VPWR _10394_/Y sky130_fd_sc_hd__inv_2
X_12133_ _12042_/A _12132_/X _12042_/A _12132_/X VGND VGND VPWR VPWR _12135_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12064_ _12014_/Y _12062_/X _12063_/Y VGND VGND VPWR VPWR _12064_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11015_ _13548_/A VGND VGND VPWR VPWR _12850_/A sky130_fd_sc_hd__buf_1
XFILLER_2_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15823_ _16125_/A _15823_/B VGND VGND VPWR VPWR _15834_/B sky130_fd_sc_hd__or2_1
X_15754_ _15674_/X _15753_/Y _15674_/X _15753_/Y VGND VGND VPWR VPWR _15807_/B sky130_fd_sc_hd__a2bb2o_1
X_14705_ _14731_/A _14731_/B VGND VGND VPWR VPWR _14796_/A sky130_fd_sc_hd__and2_1
X_12966_ _13703_/A VGND VGND VPWR VPWR _14592_/A sky130_fd_sc_hd__inv_2
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15685_ _15685_/A _15685_/B VGND VGND VPWR VPWR _15685_/Y sky130_fd_sc_hd__nand2_1
X_12897_ _12844_/A _12844_/B _12844_/Y VGND VGND VPWR VPWR _12897_/Y sky130_fd_sc_hd__o21ai_1
X_11917_ _11985_/A VGND VGND VPWR VPWR _12775_/A sky130_fd_sc_hd__buf_1
XFILLER_33_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14576_/A _14576_/B _14576_/Y VGND VGND VPWR VPWR _14636_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11848_ _11848_/A VGND VGND VPWR VPWR _11848_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14567_ _15272_/A _14574_/B VGND VGND VPWR VPWR _14567_/Y sky130_fd_sc_hd__nor2_1
X_16306_ _16253_/A _16320_/A _16253_/Y VGND VGND VPWR VPWR _16306_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11779_ _11728_/B _11778_/Y _11728_/B _11778_/Y VGND VGND VPWR VPWR _11780_/B sky130_fd_sc_hd__o2bb2a_1
X_13518_ _10476_/X _13485_/X _10476_/X _13485_/X VGND VGND VPWR VPWR _13519_/B sky130_fd_sc_hd__o2bb2a_1
X_14498_ _14461_/A _14461_/B _14461_/Y VGND VGND VPWR VPWR _14498_/Y sky130_fd_sc_hd__o21ai_1
X_16237_ _15786_/Y _16236_/X _15786_/Y _16236_/X VGND VGND VPWR VPWR _16238_/B sky130_fd_sc_hd__a2bb2oi_1
X_13449_ _13378_/Y _13447_/X _13448_/Y VGND VGND VPWR VPWR _13449_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16168_ _16192_/A _16168_/B VGND VGND VPWR VPWR _16266_/B sky130_fd_sc_hd__or2_1
XFILLER_126_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15119_ _15119_/A _15119_/B VGND VGND VPWR VPWR _15119_/Y sky130_fd_sc_hd__nand2_1
X_16099_ _16099_/A _16099_/B VGND VGND VPWR VPWR _16099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08990_ _09478_/B _08989_/Y _08514_/Y _08695_/Y VGND VGND VPWR VPWR _08990_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09611_ _09509_/X _09610_/X _09509_/X _09610_/X VGND VGND VPWR VPWR _09977_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09542_ _09629_/B VGND VGND VPWR VPWR _09628_/B sky130_fd_sc_hd__inv_2
X_09473_ _09451_/Y _09471_/X _09472_/X VGND VGND VPWR VPWR _09473_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08424_ _08424_/A VGND VGND VPWR VPWR _08424_/Y sky130_fd_sc_hd__inv_2
X_08355_ _08355_/A VGND VGND VPWR VPWR _08355_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08286_ input28/X _08352_/B _08353_/A _08355_/A VGND VGND VPWR VPWR _08349_/A sky130_fd_sc_hd__o22a_1
XFILLER_118_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09809_ _08844_/A _09230_/A _09459_/Y _09826_/A VGND VGND VPWR VPWR _09809_/X sky130_fd_sc_hd__o22a_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12820_ _12765_/A _12765_/B _12765_/Y VGND VGND VPWR VPWR _12820_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12700_/A _12700_/B _12700_/Y VGND VGND VPWR VPWR _12751_/X sky130_fd_sc_hd__a21o_1
X_15470_ _15470_/A _15470_/B VGND VGND VPWR VPWR _15470_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11696_/X _11701_/Y _11696_/X _11701_/Y VGND VGND VPWR VPWR _11702_/Y sky130_fd_sc_hd__a2bb2oi_1
X_12682_ _12682_/A _12682_/B VGND VGND VPWR VPWR _12682_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14421_ _14421_/A _14421_/B VGND VGND VPWR VPWR _14421_/Y sky130_fd_sc_hd__nor2_1
X_11633_ _11631_/Y _11632_/Y _11540_/Y VGND VGND VPWR VPWR _11633_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14352_ _13415_/Y _14351_/X _13415_/Y _14351_/X VGND VGND VPWR VPWR _14353_/B sky130_fd_sc_hd__a2bb2oi_1
X_11564_ _12407_/A _11564_/B VGND VGND VPWR VPWR _11564_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14283_ _14286_/A _15908_/A VGND VGND VPWR VPWR _14399_/A sky130_fd_sc_hd__and2_1
X_13303_ _14771_/A _13303_/B VGND VGND VPWR VPWR _13303_/Y sky130_fd_sc_hd__nand2_1
X_11495_ _09997_/B _11494_/X _09997_/B _11494_/X VGND VGND VPWR VPWR _11496_/B sky130_fd_sc_hd__o2bb2a_1
X_10515_ _09829_/A _09829_/B _09830_/A VGND VGND VPWR VPWR _10515_/Y sky130_fd_sc_hd__o21ai_1
X_16022_ _16032_/A _16032_/B VGND VGND VPWR VPWR _16022_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13234_ _13197_/X _13233_/Y _13197_/X _13233_/Y VGND VGND VPWR VPWR _13294_/B sky130_fd_sc_hd__a2bb2o_1
X_10446_ _10446_/A VGND VGND VPWR VPWR _10957_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13165_ _13192_/A _13192_/B VGND VGND VPWR VPWR _13165_/Y sky130_fd_sc_hd__nor2_1
X_10377_ _10377_/A VGND VGND VPWR VPWR _10377_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12116_ _13910_/A _12147_/B VGND VGND VPWR VPWR _12213_/A sky130_fd_sc_hd__and2_1
X_13096_ _13096_/A VGND VGND VPWR VPWR _13096_/X sky130_fd_sc_hd__buf_1
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12047_ _12047_/A _12047_/B VGND VGND VPWR VPWR _12047_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15806_ _15802_/Y _16207_/A _15805_/Y VGND VGND VPWR VPWR _16197_/A sky130_fd_sc_hd__o21ai_2
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13998_ _13998_/A VGND VGND VPWR VPWR _13998_/Y sky130_fd_sc_hd__inv_2
X_15737_ _16112_/A _15813_/B VGND VGND VPWR VPWR _15737_/Y sky130_fd_sc_hd__nor2_1
X_12949_ _12864_/X _12948_/X _12864_/X _12948_/X VGND VGND VPWR VPWR _12951_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15668_ _15785_/A _15666_/X _15667_/X VGND VGND VPWR VPWR _15668_/Y sky130_fd_sc_hd__o21ai_1
X_14619_ _14619_/A VGND VGND VPWR VPWR _15341_/A sky130_fd_sc_hd__buf_1
XFILLER_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15599_ _15681_/A _15681_/B VGND VGND VPWR VPWR _15599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08973_ _08907_/X _08971_/X _11385_/B VGND VGND VPWR VPWR _08973_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09525_ _09525_/A _09525_/B VGND VGND VPWR VPWR _09526_/A sky130_fd_sc_hd__or2_1
XFILLER_52_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09456_ _09456_/A _09456_/B VGND VGND VPWR VPWR _09456_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08407_ _09006_/A _08403_/Y _09459_/A VGND VGND VPWR VPWR _08407_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09387_ _09430_/B _09371_/B _09371_/X _11474_/A VGND VGND VPWR VPWR _11576_/A sky130_fd_sc_hd__a22o_1
X_08338_ _08338_/A VGND VGND VPWR VPWR _08338_/Y sky130_fd_sc_hd__inv_2
X_08269_ _08269_/A input12/X VGND VGND VPWR VPWR _08353_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10300_ _09717_/A _09113_/B _09113_/Y VGND VGND VPWR VPWR _10300_/X sky130_fd_sc_hd__o21a_1
X_11280_ _11583_/A _11280_/B VGND VGND VPWR VPWR _12290_/A sky130_fd_sc_hd__or2_2
XFILLER_118_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10231_ _10231_/A VGND VGND VPWR VPWR _10231_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10162_ _08810_/B _10127_/B _10128_/B VGND VGND VPWR VPWR _10163_/B sky130_fd_sc_hd__a21bo_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14970_ _14935_/X _14949_/A _14948_/X VGND VGND VPWR VPWR _14970_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10093_ _10055_/A _10055_/B _10055_/X VGND VGND VPWR VPWR _10094_/A sky130_fd_sc_hd__a21bo_1
X_13921_ _15404_/A _13946_/B VGND VGND VPWR VPWR _13921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13852_ _14615_/A _13852_/B VGND VGND VPWR VPWR _13852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13783_ _13713_/A _13713_/B _13782_/Y _13710_/X VGND VGND VPWR VPWR _13783_/X sky130_fd_sc_hd__o22a_1
X_12803_ _12776_/X _12802_/Y _12776_/X _12802_/Y VGND VGND VPWR VPWR _12852_/B sky130_fd_sc_hd__a2bb2o_1
X_15522_ _15464_/A _15464_/B _15464_/Y VGND VGND VPWR VPWR _15522_/Y sky130_fd_sc_hd__o21ai_1
X_10995_ _12160_/A _11115_/B VGND VGND VPWR VPWR _10995_/Y sky130_fd_sc_hd__nand2_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12734_ _12716_/X _12733_/X _12716_/X _12733_/X VGND VGND VPWR VPWR _12779_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15453_ _15453_/A _15408_/X VGND VGND VPWR VPWR _15453_/X sky130_fd_sc_hd__or2b_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _10673_/Y _12664_/Y _10564_/Y VGND VGND VPWR VPWR _12666_/A sky130_fd_sc_hd__o21ai_1
XFILLER_15_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14404_ _14297_/Y _14402_/X _14403_/Y VGND VGND VPWR VPWR _14404_/X sky130_fd_sc_hd__o21a_1
X_12596_ _14901_/A VGND VGND VPWR VPWR _14906_/A sky130_fd_sc_hd__buf_1
X_15384_ _15384_/A _15335_/X VGND VGND VPWR VPWR _15384_/X sky130_fd_sc_hd__or2b_1
X_11616_ _11616_/A _11616_/B VGND VGND VPWR VPWR _11616_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14335_ _14335_/A _14335_/B VGND VGND VPWR VPWR _15956_/A sky130_fd_sc_hd__or2_1
X_11547_ _12953_/A _11643_/B _11546_/Y VGND VGND VPWR VPWR _11547_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16005_ _16005_/A _15960_/X VGND VGND VPWR VPWR _16005_/X sky130_fd_sc_hd__or2b_1
X_14266_ _15866_/A _14266_/B VGND VGND VPWR VPWR _14266_/Y sky130_fd_sc_hd__nand2_1
X_11478_ _13873_/A VGND VGND VPWR VPWR _15107_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14197_ _12628_/X _14196_/X _12628_/X _14196_/X VGND VGND VPWR VPWR _14269_/B sky130_fd_sc_hd__a2bb2o_1
X_13217_ _14754_/A VGND VGND VPWR VPWR _14771_/A sky130_fd_sc_hd__buf_1
X_10429_ _10429_/A VGND VGND VPWR VPWR _11791_/A sky130_fd_sc_hd__buf_1
XFILLER_124_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13148_ _15240_/A _13121_/B _13121_/Y VGND VGND VPWR VPWR _13148_/Y sky130_fd_sc_hd__o21ai_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _13763_/A VGND VGND VPWR VPWR _15258_/A sky130_fd_sc_hd__buf_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09310_ _10252_/A _09310_/B VGND VGND VPWR VPWR _09310_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09241_ _08623_/A _09802_/A _09224_/Y _09240_/Y VGND VGND VPWR VPWR _09241_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09172_ _09754_/A VGND VGND VPWR VPWR _09430_/A sky130_fd_sc_hd__buf_1
XFILLER_119_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08956_ _08954_/Y _08955_/Y _08954_/Y _08955_/Y VGND VGND VPWR VPWR _08960_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08887_ _08687_/X _08886_/Y _08687_/X _08886_/Y VGND VGND VPWR VPWR _08978_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09508_ _09500_/A _09500_/B _09500_/Y _09507_/X VGND VGND VPWR VPWR _09508_/X sky130_fd_sc_hd__o2bb2a_1
X_10780_ _12066_/A VGND VGND VPWR VPWR _13058_/A sky130_fd_sc_hd__buf_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09439_ _09431_/A _09431_/B _09431_/X _09438_/X VGND VGND VPWR VPWR _09439_/X sky130_fd_sc_hd__a22o_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _12449_/Y _12366_/X _12387_/Y VGND VGND VPWR VPWR _12450_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11401_ _08952_/A _08952_/B _08952_/Y VGND VGND VPWR VPWR _11401_/X sky130_fd_sc_hd__o21a_1
X_14120_ _14120_/A VGND VGND VPWR VPWR _14876_/A sky130_fd_sc_hd__inv_2
X_12381_ _12417_/B _12380_/X _12417_/B _12380_/X VGND VGND VPWR VPWR _12382_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11332_ _11516_/A _12373_/A _11331_/Y VGND VGND VPWR VPWR _11332_/X sky130_fd_sc_hd__a21o_1
X_14051_ _14039_/A _14039_/B _14039_/X _14050_/X VGND VGND VPWR VPWR _14051_/X sky130_fd_sc_hd__o22a_1
X_11263_ _11263_/A VGND VGND VPWR VPWR _11263_/Y sky130_fd_sc_hd__inv_2
X_11194_ _14058_/A VGND VGND VPWR VPWR _15449_/A sky130_fd_sc_hd__buf_1
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13002_ _13002_/A VGND VGND VPWR VPWR _13002_/X sky130_fd_sc_hd__buf_1
X_10214_ _10201_/Y _10212_/X _10213_/Y VGND VGND VPWR VPWR _10309_/B sky130_fd_sc_hd__o21ai_2
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10145_ _10147_/A VGND VGND VPWR VPWR _10240_/B sky130_fd_sc_hd__buf_1
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14953_ _14953_/A _14953_/B VGND VGND VPWR VPWR _14953_/Y sky130_fd_sc_hd__nor2_1
X_10076_ _10075_/A _10075_/B _09700_/A _10075_/X VGND VGND VPWR VPWR _10076_/X sky130_fd_sc_hd__a22o_1
X_14884_ _14794_/A _14794_/B _14794_/A _14794_/B VGND VGND VPWR VPWR _14884_/X sky130_fd_sc_hd__a2bb2o_1
X_13904_ _13853_/X _13903_/Y _13853_/X _13903_/Y VGND VGND VPWR VPWR _13954_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13835_ _13753_/A _13753_/B _13753_/Y VGND VGND VPWR VPWR _13835_/Y sky130_fd_sc_hd__a21oi_1
X_13766_ _13816_/A _13764_/X _13765_/X VGND VGND VPWR VPWR _13766_/X sky130_fd_sc_hd__o21a_1
X_10978_ _10978_/A VGND VGND VPWR VPWR _10978_/Y sky130_fd_sc_hd__inv_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15505_ _15480_/X _15504_/X _15480_/X _15504_/X VGND VGND VPWR VPWR _15542_/B sky130_fd_sc_hd__a2bb2o_1
X_13697_ _13697_/A _13697_/B VGND VGND VPWR VPWR _13697_/X sky130_fd_sc_hd__or2_1
X_12717_ _12688_/A _12688_/B _12688_/Y _12716_/X VGND VGND VPWR VPWR _12717_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12648_ _12648_/A _12648_/B VGND VGND VPWR VPWR _12650_/B sky130_fd_sc_hd__or2_1
X_15436_ _15419_/X _15435_/X _15419_/X _15435_/X VGND VGND VPWR VPWR _15437_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12579_ _12574_/Y _12578_/Y _12574_/A _12578_/A _11706_/A VGND VGND VPWR VPWR _12621_/A
+ sky130_fd_sc_hd__o221a_1
X_15367_ _15346_/X _15366_/X _15346_/X _15366_/X VGND VGND VPWR VPWR _15414_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14318_ _15962_/A _14392_/B VGND VGND VPWR VPWR _15597_/A sky130_fd_sc_hd__and2_1
X_15298_ _15281_/X _15297_/Y _15281_/X _15297_/Y VGND VGND VPWR VPWR _15349_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14249_ _14372_/B _14249_/B VGND VGND VPWR VPWR _15885_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08810_ _10015_/A _08810_/B VGND VGND VPWR VPWR _08810_/Y sky130_fd_sc_hd__nor2_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09169_/A _09749_/X _09750_/Y _09789_/X VGND VGND VPWR VPWR _09793_/A sky130_fd_sc_hd__o22a_1
XFILLER_97_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08741_ _08710_/Y _08739_/Y _08740_/X VGND VGND VPWR VPWR _08742_/A sky130_fd_sc_hd__o21ai_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08672_ _09680_/A VGND VGND VPWR VPWR _10098_/A sky130_fd_sc_hd__inv_2
XFILLER_54_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09224_ _09224_/A VGND VGND VPWR VPWR _09224_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09155_ _09527_/B _09155_/B VGND VGND VPWR VPWR _09156_/B sky130_fd_sc_hd__or2_1
X_09086_ _09769_/A VGND VGND VPWR VPWR _09424_/A sky130_fd_sc_hd__buf_1
XFILLER_123_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09988_ _09968_/Y _09986_/Y _09987_/Y VGND VGND VPWR VPWR _09990_/B sky130_fd_sc_hd__o21ai_2
X_08939_ _08942_/A _08942_/B VGND VGND VPWR VPWR _08939_/Y sky130_fd_sc_hd__nor2_1
X_11950_ _11897_/A _11949_/Y _11897_/A _11949_/Y VGND VGND VPWR VPWR _11968_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10901_ _10901_/A _10766_/X VGND VGND VPWR VPWR _10901_/X sky130_fd_sc_hd__or2b_1
XFILLER_57_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11881_ _11836_/X _11880_/Y _11836_/X _11880_/Y VGND VGND VPWR VPWR _11895_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13620_ _15140_/A _13606_/B _13606_/Y _13619_/X VGND VGND VPWR VPWR _13620_/X sky130_fd_sc_hd__o2bb2a_1
X_10832_ _13510_/A _10953_/B _13510_/A _10953_/B VGND VGND VPWR VPWR _10832_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10763_ _15212_/A _12041_/A VGND VGND VPWR VPWR _13006_/A sky130_fd_sc_hd__or2_1
X_13551_ _13536_/X _13550_/Y _13536_/X _13550_/Y VGND VGND VPWR VPWR _13552_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16270_ _16270_/A _16270_/B VGND VGND VPWR VPWR _16270_/Y sky130_fd_sc_hd__nand2_1
X_12502_ _12409_/A _12409_/B _12409_/Y _12501_/X VGND VGND VPWR VPWR _12639_/B sky130_fd_sc_hd__o211a_1
XFILLER_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15221_ _15202_/A _15202_/B _15202_/Y _15220_/X VGND VGND VPWR VPWR _15221_/X sky130_fd_sc_hd__a2bb2o_1
X_13482_ _11731_/A _10294_/Y _10335_/Y _13481_/Y VGND VGND VPWR VPWR _13482_/X sky130_fd_sc_hd__o22a_1
X_10694_ _13513_/A _10801_/B _13513_/A _10801_/B VGND VGND VPWR VPWR _10694_/X sky130_fd_sc_hd__a2bb2o_1
X_12433_ _13495_/A _12432_/B _12432_/Y VGND VGND VPWR VPWR _12437_/A sky130_fd_sc_hd__a21oi_1
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12364_ _12362_/Y _12363_/Y _12284_/Y VGND VGND VPWR VPWR _12364_/X sky130_fd_sc_hd__o21a_1
X_15152_ _15131_/A _15131_/B _15131_/Y _15151_/X VGND VGND VPWR VPWR _15152_/X sky130_fd_sc_hd__a2bb2o_1
X_14103_ _14103_/A _14106_/B VGND VGND VPWR VPWR _14103_/Y sky130_fd_sc_hd__nor2_1
X_15083_ _15027_/X _15082_/X _15027_/X _15082_/X VGND VGND VPWR VPWR _15084_/B sky130_fd_sc_hd__a2bb2o_1
X_11315_ _11314_/Y _11141_/X _11150_/Y VGND VGND VPWR VPWR _11315_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14034_ _15402_/A _13944_/B _13944_/Y VGND VGND VPWR VPWR _14034_/Y sky130_fd_sc_hd__o21ai_1
X_12295_ _12295_/A _12294_/X VGND VGND VPWR VPWR _12295_/X sky130_fd_sc_hd__or2b_1
X_11246_ _11246_/A _11072_/X VGND VGND VPWR VPWR _11246_/X sky130_fd_sc_hd__or2b_1
X_11177_ _11177_/A _11176_/X VGND VGND VPWR VPWR _11177_/X sky130_fd_sc_hd__or2b_1
X_15985_ _15984_/Y _15979_/X _15976_/Y VGND VGND VPWR VPWR _15985_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10128_ _10128_/A _10128_/B VGND VGND VPWR VPWR _10129_/B sky130_fd_sc_hd__or2_1
X_14936_ _12785_/A _12382_/B _12382_/Y _14839_/X VGND VGND VPWR VPWR _14936_/X sky130_fd_sc_hd__o2bb2a_1
X_10059_ _10059_/A _10059_/B VGND VGND VPWR VPWR _10059_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14867_ _15550_/A _14926_/B VGND VGND VPWR VPWR _14867_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14798_ _14798_/A _14798_/B VGND VGND VPWR VPWR _14798_/X sky130_fd_sc_hd__and2_1
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13818_ _14623_/A _13848_/B VGND VGND VPWR VPWR _13818_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13749_ _13686_/A _13748_/Y _13686_/A _13748_/Y VGND VGND VPWR VPWR _13757_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16468_ _16357_/A _16468_/D VGND VGND VPWR VPWR _16468_/Q sky130_fd_sc_hd__dfxtp_1
X_16399_ _16402_/B VGND VGND VPWR VPWR _16399_/Y sky130_fd_sc_hd__inv_2
X_15419_ _15438_/A _15417_/X _15418_/X VGND VGND VPWR VPWR _15419_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09911_ _09911_/A _09910_/Y VGND VGND VPWR VPWR _09913_/B sky130_fd_sc_hd__or2b_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09842_ _09843_/A _09843_/B VGND VGND VPWR VPWR _10491_/A sky130_fd_sc_hd__and2_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A _09773_/B VGND VGND VPWR VPWR _09773_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08724_ _09228_/A _09458_/B VGND VGND VPWR VPWR _08724_/X sky130_fd_sc_hd__or2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08655_ _09799_/A VGND VGND VPWR VPWR _09684_/A sky130_fd_sc_hd__inv_2
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08586_ _08586_/A VGND VGND VPWR VPWR _08586_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09207_ _14012_/A VGND VGND VPWR VPWR _14062_/A sky130_fd_sc_hd__buf_1
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09138_ _09436_/A _09141_/B VGND VGND VPWR VPWR _09138_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11100_ _13713_/A VGND VGND VPWR VPWR _12856_/A sky130_fd_sc_hd__buf_1
X_09069_ _09069_/A _09069_/B VGND VGND VPWR VPWR _09070_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12080_ _12080_/A _12080_/B VGND VGND VPWR VPWR _12080_/X sky130_fd_sc_hd__or2_1
XFILLER_1_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11031_ _15072_/A VGND VGND VPWR VPWR _13914_/A sky130_fd_sc_hd__buf_1
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15770_ _15770_/A VGND VGND VPWR VPWR _15770_/Y sky130_fd_sc_hd__inv_2
X_12982_ _13695_/A VGND VGND VPWR VPWR _14485_/A sky130_fd_sc_hd__inv_2
X_14721_ _14722_/A _14722_/B VGND VGND VPWR VPWR _14721_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11933_ _11933_/A _11981_/B VGND VGND VPWR VPWR _11933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14652_ _15337_/A _14652_/B VGND VGND VPWR VPWR _14652_/Y sky130_fd_sc_hd__nand2_1
X_11864_ _11913_/B _11863_/Y _11913_/B _11863_/Y VGND VGND VPWR VPWR _11911_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13603_ _13606_/A VGND VGND VPWR VPWR _15140_/A sky130_fd_sc_hd__buf_1
X_10815_ _10966_/A _10815_/B VGND VGND VPWR VPWR _10816_/A sky130_fd_sc_hd__or2_1
X_16322_ _16322_/A _16322_/B VGND VGND VPWR VPWR _16322_/Y sky130_fd_sc_hd__nand2_1
X_14583_ _14551_/Y _14581_/X _14582_/Y VGND VGND VPWR VPWR _14583_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11795_ _13568_/A _11780_/B _11780_/X _11794_/X VGND VGND VPWR VPWR _11795_/X sky130_fd_sc_hd__o22a_1
XFILLER_41_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10746_ _10631_/A _10745_/Y _10631_/A _10745_/Y VGND VGND VPWR VPWR _10747_/B sky130_fd_sc_hd__a2bb2o_1
X_13534_ _15032_/A _13525_/B _13525_/Y _13533_/X VGND VGND VPWR VPWR _13534_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16253_ _16253_/A _16253_/B VGND VGND VPWR VPWR _16253_/Y sky130_fd_sc_hd__nand2_1
X_13465_ _13462_/Y _13464_/X _13462_/Y _13464_/X VGND VGND VPWR VPWR _13465_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10677_ _10966_/A _10677_/B VGND VGND VPWR VPWR _10678_/A sky130_fd_sc_hd__or2_1
X_16184_ _16192_/A _16184_/B VGND VGND VPWR VPWR _16262_/B sky130_fd_sc_hd__or2_1
X_15204_ _15149_/X _15203_/Y _15149_/X _15203_/Y VGND VGND VPWR VPWR _15205_/B sky130_fd_sc_hd__a2bb2o_1
X_12416_ _12416_/A VGND VGND VPWR VPWR _12682_/A sky130_fd_sc_hd__buf_1
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13396_ _13396_/A VGND VGND VPWR VPWR _14098_/A sky130_fd_sc_hd__inv_2
XFILLER_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15135_ _15078_/A _15078_/B _15078_/Y VGND VGND VPWR VPWR _15135_/Y sky130_fd_sc_hd__o21ai_1
X_12347_ _11449_/A _12215_/B _12215_/Y VGND VGND VPWR VPWR _12347_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15066_ _15066_/A _15066_/B VGND VGND VPWR VPWR _15066_/Y sky130_fd_sc_hd__nand2_1
X_12278_ _12369_/B _12277_/Y _12369_/B _12277_/Y VGND VGND VPWR VPWR _12367_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14017_ _13953_/X _14016_/Y _13953_/X _14016_/Y VGND VGND VPWR VPWR _14058_/B sky130_fd_sc_hd__a2bb2o_1
X_11229_ _11080_/X _11228_/X _11080_/X _11228_/X VGND VGND VPWR VPWR _11230_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15968_ _15905_/X _15967_/Y _15905_/X _15967_/Y VGND VGND VPWR VPWR _15968_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15899_ _15865_/Y _15897_/X _15898_/Y VGND VGND VPWR VPWR _15899_/X sky130_fd_sc_hd__o21a_1
X_14919_ _14883_/Y _14917_/X _14918_/Y VGND VGND VPWR VPWR _14919_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08440_ _08440_/A VGND VGND VPWR VPWR _08440_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08371_ input15/X _08260_/B _08337_/B _08424_/A VGND VGND VPWR VPWR _08429_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09825_ _09818_/A _09818_/B _09819_/B VGND VGND VPWR VPWR _09838_/A sky130_fd_sc_hd__a21bo_1
XFILLER_101_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09756_ _10085_/A VGND VGND VPWR VPWR _09995_/B sky130_fd_sc_hd__buf_1
XFILLER_100_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08707_ _09448_/B VGND VGND VPWR VPWR _08755_/A sky130_fd_sc_hd__inv_2
X_09687_ _09687_/A _09687_/B VGND VGND VPWR VPWR _09690_/B sky130_fd_sc_hd__or2_1
XFILLER_27_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08483_/X _08388_/A _08483_/X _08388_/A VGND VGND VPWR VPWR _08639_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _09453_/B VGND VGND VPWR VPWR _08713_/B sky130_fd_sc_hd__inv_2
X_11580_ _11555_/A _11481_/X _11554_/X VGND VGND VPWR VPWR _11580_/X sky130_fd_sc_hd__o21a_1
X_10600_ _10735_/A _10635_/B VGND VGND VPWR VPWR _10600_/Y sky130_fd_sc_hd__nor2_1
X_10531_ _11841_/A _10531_/B VGND VGND VPWR VPWR _10531_/Y sky130_fd_sc_hd__nand2_1
X_13250_ _14731_/A _13285_/B VGND VGND VPWR VPWR _13250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12201_ _12201_/A _12200_/X VGND VGND VPWR VPWR _12201_/X sky130_fd_sc_hd__or2b_1
XFILLER_89_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10462_ _10462_/A VGND VGND VPWR VPWR _10462_/Y sky130_fd_sc_hd__inv_2
X_13181_ _13096_/X _13180_/Y _13096_/A _13180_/Y VGND VGND VPWR VPWR _13182_/B sky130_fd_sc_hd__a2bb2o_1
X_10393_ _10245_/A _09307_/B _09307_/Y VGND VGND VPWR VPWR _10394_/A sky130_fd_sc_hd__o21ai_1
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12132_ _12047_/A _12047_/B _12047_/Y VGND VGND VPWR VPWR _12132_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12063_ _12063_/A _12063_/B VGND VGND VPWR VPWR _12063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11014_ _11014_/A VGND VGND VPWR VPWR _13548_/A sky130_fd_sc_hd__buf_1
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15822_ _15712_/X _15820_/X _16142_/B VGND VGND VPWR VPWR _15822_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15753_ _15675_/A _15675_/B _15675_/Y VGND VGND VPWR VPWR _15753_/Y sky130_fd_sc_hd__o21ai_1
X_12965_ _14669_/A _13030_/B VGND VGND VPWR VPWR _13050_/A sky130_fd_sc_hd__and2_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14704_ _14653_/X _14703_/Y _14653_/X _14703_/Y VGND VGND VPWR VPWR _14731_/B sky130_fd_sc_hd__a2bb2o_1
X_11916_ _11916_/A VGND VGND VPWR VPWR _11985_/A sky130_fd_sc_hd__inv_2
XFILLER_45_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15684_ _15592_/Y _15682_/X _15683_/Y VGND VGND VPWR VPWR _15684_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12896_ _12930_/A VGND VGND VPWR VPWR _14465_/A sky130_fd_sc_hd__buf_1
XFILLER_45_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14635_/A VGND VGND VPWR VPWR _15333_/A sky130_fd_sc_hd__buf_1
XFILLER_60_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11847_ _11847_/A _11847_/B VGND VGND VPWR VPWR _11847_/X sky130_fd_sc_hd__or2_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14509_/X _14565_/X _14509_/X _14565_/X VGND VGND VPWR VPWR _14574_/B sky130_fd_sc_hd__a2bb2o_1
X_11778_ _12765_/A _11777_/B _11777_/Y VGND VGND VPWR VPWR _11778_/Y sky130_fd_sc_hd__a21oi_1
X_16305_ _16322_/A _16322_/B VGND VGND VPWR VPWR _16305_/Y sky130_fd_sc_hd__nor2_1
X_10729_ _11970_/A _10729_/B VGND VGND VPWR VPWR _10729_/Y sky130_fd_sc_hd__nand2_1
X_13517_ _13519_/A VGND VGND VPWR VPWR _15036_/A sky130_fd_sc_hd__buf_1
XFILLER_41_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16236_ _16089_/A _15788_/B _15788_/Y VGND VGND VPWR VPWR _16236_/X sky130_fd_sc_hd__o21a_1
X_14497_ _14497_/A VGND VGND VPWR VPWR _15208_/A sky130_fd_sc_hd__buf_1
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13448_ _13448_/A _13448_/B VGND VGND VPWR VPWR _13448_/Y sky130_fd_sc_hd__nand2_1
X_16167_ _15814_/X _16166_/X _15814_/X _16166_/X VGND VGND VPWR VPWR _16168_/B sky130_fd_sc_hd__a2bb2o_1
X_13379_ _13379_/A _13371_/X VGND VGND VPWR VPWR _13379_/X sky130_fd_sc_hd__or2b_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16098_ _16033_/X _16097_/Y _16033_/X _16097_/Y VGND VGND VPWR VPWR _16098_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15118_ _15096_/X _15117_/Y _15096_/X _15117_/Y VGND VGND VPWR VPWR _15119_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15049_ _12274_/X _15048_/X _12274_/X _15048_/X VGND VGND VPWR VPWR _15051_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09610_ _09496_/A _09496_/B _09496_/Y VGND VGND VPWR VPWR _09610_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09541_ _09541_/A _09541_/B VGND VGND VPWR VPWR _09629_/B sky130_fd_sc_hd__or2_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09472_ _10011_/A _09472_/B VGND VGND VPWR VPWR _09472_/X sky130_fd_sc_hd__or2_1
X_08423_ _09217_/B _08417_/Y _09250_/A VGND VGND VPWR VPWR _08423_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08354_ _08354_/A VGND VGND VPWR VPWR _08354_/Y sky130_fd_sc_hd__inv_2
X_08285_ input27/X _08363_/B _08364_/A _08384_/A VGND VGND VPWR VPWR _08355_/A sky130_fd_sc_hd__o22a_1
XFILLER_118_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09808_ _09808_/A VGND VGND VPWR VPWR _09826_/A sky130_fd_sc_hd__inv_2
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09739_ _09739_/A _09739_/B VGND VGND VPWR VPWR _09742_/A sky130_fd_sc_hd__or2_1
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12750_ _12769_/A _12769_/B VGND VGND VPWR VPWR _12750_/Y sky130_fd_sc_hd__nor2_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11701_ _11697_/X _11700_/X _11697_/X _11700_/X VGND VGND VPWR VPWR _11701_/Y sky130_fd_sc_hd__a2bb2oi_1
X_12681_ _11530_/A _12676_/A _11530_/Y _12676_/Y VGND VGND VPWR VPWR _12682_/B sky130_fd_sc_hd__o22a_1
XFILLER_91_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _11814_/Y _14419_/X _11814_/Y _14419_/X VGND VGND VPWR VPWR _14421_/B sky130_fd_sc_hd__o2bb2a_1
X_11632_ _11632_/A VGND VGND VPWR VPWR _11632_/Y sky130_fd_sc_hd__inv_2
X_14351_ _13413_/X _14351_/B VGND VGND VPWR VPWR _14351_/X sky130_fd_sc_hd__and2b_1
X_11563_ _11466_/X _11562_/Y _11466_/X _11562_/Y VGND VGND VPWR VPWR _11564_/B sky130_fd_sc_hd__a2bb2o_1
X_13302_ _13302_/A VGND VGND VPWR VPWR _13302_/Y sky130_fd_sc_hd__inv_2
X_14282_ _14282_/A _14282_/B VGND VGND VPWR VPWR _15908_/A sky130_fd_sc_hd__or2_1
XFILLER_109_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10514_ _15143_/A _10525_/B VGND VGND VPWR VPWR _10514_/Y sky130_fd_sc_hd__nor2_1
X_11494_ _11494_/A _09788_/X VGND VGND VPWR VPWR _11494_/X sky130_fd_sc_hd__or2b_1
XFILLER_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16021_ _15949_/X _16020_/X _15949_/X _16020_/X VGND VGND VPWR VPWR _16032_/B sky130_fd_sc_hd__a2bb2o_1
X_13233_ _13198_/A _13198_/B _13198_/Y VGND VGND VPWR VPWR _13233_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10445_ _10445_/A VGND VGND VPWR VPWR _10445_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13164_ _13110_/X _13163_/Y _13110_/X _13163_/Y VGND VGND VPWR VPWR _13192_/B sky130_fd_sc_hd__a2bb2o_1
X_12115_ _12058_/X _12114_/Y _12058_/X _12114_/Y VGND VGND VPWR VPWR _12147_/B sky130_fd_sc_hd__a2bb2o_1
X_10376_ _10376_/A VGND VGND VPWR VPWR _10376_/Y sky130_fd_sc_hd__inv_2
X_13095_ _14564_/A _13103_/B VGND VGND VPWR VPWR _13095_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12046_ _13833_/A _12047_/B VGND VGND VPWR VPWR _12046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15805_ _16104_/A _15805_/B VGND VGND VPWR VPWR _15805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13997_ _13544_/X _13996_/Y _13544_/X _13996_/Y VGND VGND VPWR VPWR _13997_/X sky130_fd_sc_hd__a2bb2o_1
X_15736_ _15680_/X _15735_/Y _15680_/X _15735_/Y VGND VGND VPWR VPWR _15813_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12948_ _12867_/Y _12945_/X _12947_/Y VGND VGND VPWR VPWR _12948_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15667_ _15667_/A _15667_/B VGND VGND VPWR VPWR _15667_/X sky130_fd_sc_hd__or2_1
X_12879_ _14600_/A _12940_/B VGND VGND VPWR VPWR _12879_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14618_ _15343_/A _14658_/B VGND VGND VPWR VPWR _14618_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15598_ _14391_/X _15597_/X _14391_/X _15597_/X VGND VGND VPWR VPWR _15681_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14549_ _14549_/A _14518_/X VGND VGND VPWR VPWR _14549_/X sky130_fd_sc_hd__or2b_1
X_16219_ _16217_/A _16218_/A _16217_/Y _16218_/Y _15832_/A VGND VGND VPWR VPWR _16253_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08972_ _08972_/A _08972_/B VGND VGND VPWR VPWR _11385_/B sky130_fd_sc_hd__or2_1
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09524_ _09561_/A _09561_/B VGND VGND VPWR VPWR _09567_/A sky130_fd_sc_hd__nor2_1
X_09455_ _09494_/A _09455_/B VGND VGND VPWR VPWR _09455_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08406_ _08944_/A VGND VGND VPWR VPWR _09459_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09386_ _09431_/B _09377_/B _09377_/X _11269_/A VGND VGND VPWR VPWR _11474_/A sky130_fd_sc_hd__a22o_1
X_08337_ _08337_/A _08337_/B VGND VGND VPWR VPWR _08338_/A sky130_fd_sc_hd__or2_1
XFILLER_20_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08268_ input28/X VGND VGND VPWR VPWR _08269_/A sky130_fd_sc_hd__inv_2
XFILLER_106_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10230_ _10230_/A _10230_/B VGND VGND VPWR VPWR _10231_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10161_ _10163_/A VGND VGND VPWR VPWR _10244_/B sky130_fd_sc_hd__buf_1
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10092_ _10007_/X _10091_/X _10007_/X _10091_/X VGND VGND VPWR VPWR _10215_/A sky130_fd_sc_hd__a2bb2o_4
X_13920_ _13845_/X _13919_/Y _13845_/X _13919_/Y VGND VGND VPWR VPWR _13946_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13851_ _13815_/Y _13849_/X _13850_/Y VGND VGND VPWR VPWR _13851_/X sky130_fd_sc_hd__o21a_1
X_10994_ _10945_/X _10993_/Y _10945_/X _10993_/Y VGND VGND VPWR VPWR _11115_/B sky130_fd_sc_hd__a2bb2o_1
X_13782_ _13782_/A VGND VGND VPWR VPWR _13782_/Y sky130_fd_sc_hd__inv_2
X_12802_ _12777_/A _12777_/B _12777_/Y VGND VGND VPWR VPWR _12802_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15521_ _15524_/A _15524_/B VGND VGND VPWR VPWR _15521_/Y sky130_fd_sc_hd__nor2_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _12688_/A _12688_/B _12688_/Y VGND VGND VPWR VPWR _12733_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15452_ _15452_/A _15452_/B VGND VGND VPWR VPWR _15452_/X sky130_fd_sc_hd__and2_1
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14403_ _15972_/A _14403_/B VGND VGND VPWR VPWR _14403_/Y sky130_fd_sc_hd__nand2_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12664_/A VGND VGND VPWR VPWR _12664_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12595_ _14084_/A VGND VGND VPWR VPWR _14901_/A sky130_fd_sc_hd__buf_1
X_15383_ _15404_/A _15404_/B VGND VGND VPWR VPWR _15459_/A sky130_fd_sc_hd__and2_1
X_11615_ _11615_/A VGND VGND VPWR VPWR _11616_/B sky130_fd_sc_hd__inv_2
X_14334_ _13430_/Y _14333_/X _13430_/Y _14333_/X VGND VGND VPWR VPWR _14335_/B sky130_fd_sc_hd__a2bb2oi_1
X_11546_ _12953_/A _11643_/B VGND VGND VPWR VPWR _11546_/Y sky130_fd_sc_hd__nand2_1
X_14265_ _14265_/A VGND VGND VPWR VPWR _14265_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16004_ _16044_/A _16044_/B VGND VGND VPWR VPWR _16004_/Y sky130_fd_sc_hd__nor2_1
X_13216_ _15054_/A VGND VGND VPWR VPWR _14754_/A sky130_fd_sc_hd__inv_2
X_11477_ _13872_/A VGND VGND VPWR VPWR _13873_/A sky130_fd_sc_hd__buf_1
XFILLER_7_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14196_ _14196_/A _12629_/X VGND VGND VPWR VPWR _14196_/X sky130_fd_sc_hd__or2b_1
X_10428_ _10622_/A VGND VGND VPWR VPWR _10428_/X sky130_fd_sc_hd__buf_1
XFILLER_112_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13147_ _13204_/A _13204_/B VGND VGND VPWR VPWR _13147_/Y sky130_fd_sc_hd__nor2_1
X_10359_ _13528_/A _10328_/B _10328_/X _10358_/X VGND VGND VPWR VPWR _10359_/X sky130_fd_sc_hd__o22a_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13078_ _13078_/A VGND VGND VPWR VPWR _13763_/A sky130_fd_sc_hd__inv_2
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12029_ _11969_/X _12028_/Y _11969_/X _12028_/Y VGND VGND VPWR VPWR _12055_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15719_ _15548_/A _14924_/B _14924_/Y VGND VGND VPWR VPWR _15719_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09240_ _09458_/B _09690_/A _09227_/X _09239_/X VGND VGND VPWR VPWR _09240_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09171_ _10009_/B _09166_/B _09167_/B VGND VGND VPWR VPWR _09754_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08955_ _08955_/A VGND VGND VPWR VPWR _08955_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08886_ _08886_/A _08886_/B VGND VGND VPWR VPWR _08886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09507_ _09502_/A _09502_/B _09502_/Y _09506_/X VGND VGND VPWR VPWR _09507_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ _09432_/A _09432_/B _09432_/X _11106_/A VGND VGND VPWR VPWR _09438_/X sky130_fd_sc_hd__a22o_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09369_ _09337_/X _08873_/Y _09337_/X _08873_/Y VGND VGND VPWR VPWR _10238_/A sky130_fd_sc_hd__o2bb2a_1
X_12380_ _12380_/A _12379_/X VGND VGND VPWR VPWR _12380_/X sky130_fd_sc_hd__or2b_1
X_11400_ _11397_/Y _11399_/Y _11397_/A _11399_/A _12605_/B VGND VGND VPWR VPWR _12575_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_126_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11331_ _11516_/A _12373_/A VGND VGND VPWR VPWR _11331_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14050_ _14812_/A _14043_/B _14043_/Y _14049_/X VGND VGND VPWR VPWR _14050_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11262_ _09431_/A _09180_/B _09180_/Y VGND VGND VPWR VPWR _11263_/A sky130_fd_sc_hd__o21ai_1
XFILLER_121_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11193_ _14018_/A VGND VGND VPWR VPWR _14058_/A sky130_fd_sc_hd__buf_1
XFILLER_79_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13001_ _13001_/A VGND VGND VPWR VPWR _14505_/A sky130_fd_sc_hd__buf_1
X_10213_ _10213_/A _10213_/B VGND VGND VPWR VPWR _10213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10144_ _10118_/A _10118_/B _10119_/A VGND VGND VPWR VPWR _10147_/A sky130_fd_sc_hd__a21bo_1
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14952_ _14976_/A _14976_/B _14951_/Y VGND VGND VPWR VPWR _14952_/Y sky130_fd_sc_hd__o21ai_1
X_10075_ _10075_/A _10075_/B VGND VGND VPWR VPWR _10075_/X sky130_fd_sc_hd__or2_1
X_14883_ _15542_/A _14918_/B VGND VGND VPWR VPWR _14883_/Y sky130_fd_sc_hd__nor2_1
X_13903_ _14611_/A _13854_/B _13854_/Y VGND VGND VPWR VPWR _13903_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13834_ _13838_/A VGND VGND VPWR VPWR _14644_/A sky130_fd_sc_hd__buf_1
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13765_ _13765_/A _13765_/B VGND VGND VPWR VPWR _13765_/X sky130_fd_sc_hd__or2_1
XFILLER_50_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10977_ _12174_/A _11140_/B _10976_/Y VGND VGND VPWR VPWR _10978_/A sky130_fd_sc_hd__o21ai_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15504_ _15452_/A _15452_/B _15452_/A _15452_/B VGND VGND VPWR VPWR _15504_/X sky130_fd_sc_hd__a2bb2o_1
X_13696_ _13736_/A _13694_/X _13695_/X VGND VGND VPWR VPWR _13696_/X sky130_fd_sc_hd__o21a_1
X_12716_ _12690_/A _12690_/B _12690_/Y _12715_/X VGND VGND VPWR VPWR _12716_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12647_ _12493_/Y _12646_/X _12493_/Y _12646_/X VGND VGND VPWR VPWR _12648_/B sky130_fd_sc_hd__a2bb2oi_1
X_15435_ _15435_/A _15420_/X VGND VGND VPWR VPWR _15435_/X sky130_fd_sc_hd__or2b_1
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15366_ _15366_/A _15347_/X VGND VGND VPWR VPWR _15366_/X sky130_fd_sc_hd__or2b_1
XFILLER_129_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12578_ _12578_/A VGND VGND VPWR VPWR _12578_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14317_ _14271_/A _14316_/Y _14271_/A _14316_/Y VGND VGND VPWR VPWR _14392_/B sky130_fd_sc_hd__a2bb2o_1
X_15297_ _14746_/A _15240_/B _15240_/Y VGND VGND VPWR VPWR _15297_/Y sky130_fd_sc_hd__o21ai_1
X_11529_ _11612_/A _11612_/B _11528_/X VGND VGND VPWR VPWR _11530_/A sky130_fd_sc_hd__o21ai_1
X_14248_ _14248_/A _15838_/A VGND VGND VPWR VPWR _14249_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14179_ _12634_/X _14178_/X _12634_/X _14178_/X VGND VGND VPWR VPWR _14278_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_98_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08740_ _10010_/A _09527_/A VGND VGND VPWR VPWR _08740_/X sky130_fd_sc_hd__or2_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08671_ _08671_/A _08929_/A VGND VGND VPWR VPWR _09680_/A sky130_fd_sc_hd__or2_1
XFILLER_26_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09223_ _09547_/A _09693_/A VGND VGND VPWR VPWR _09224_/A sky130_fd_sc_hd__or2_1
XFILLER_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09154_ _09154_/A VGND VGND VPWR VPWR _09527_/B sky130_fd_sc_hd__inv_2
XFILLER_22_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09085_ _10014_/B _09075_/B _09076_/B VGND VGND VPWR VPWR _09769_/A sky130_fd_sc_hd__a21bo_1
XFILLER_122_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09987_ _09987_/A _09987_/B VGND VGND VPWR VPWR _09987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08938_ _08936_/Y _08937_/X _08936_/Y _08937_/X VGND VGND VPWR VPWR _08942_/B sky130_fd_sc_hd__a2bb2o_1
X_08869_ _08753_/Y _08868_/Y _08753_/Y _08868_/Y VGND VGND VPWR VPWR _08986_/B sky130_fd_sc_hd__o2bb2a_1
X_10900_ _12047_/A VGND VGND VPWR VPWR _13833_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11880_ _13606_/A _11837_/B _11837_/Y VGND VGND VPWR VPWR _11880_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10831_ _10810_/X _10830_/X _10810_/X _10830_/X VGND VGND VPWR VPWR _10953_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10762_ _13754_/A VGND VGND VPWR VPWR _11061_/A sky130_fd_sc_hd__inv_2
X_13550_ _15038_/A _13516_/B _13516_/Y VGND VGND VPWR VPWR _13550_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12501_ _12501_/A VGND VGND VPWR VPWR _12501_/X sky130_fd_sc_hd__clkbuf_2
X_13481_ _13481_/A VGND VGND VPWR VPWR _13481_/Y sky130_fd_sc_hd__inv_2
X_15220_ _15205_/A _15205_/B _15205_/Y _15219_/X VGND VGND VPWR VPWR _15220_/X sky130_fd_sc_hd__a2bb2o_1
X_12432_ _13495_/A _12432_/B VGND VGND VPWR VPWR _12432_/Y sky130_fd_sc_hd__nor2_1
X_10693_ _10672_/X _10692_/X _10672_/X _10692_/X VGND VGND VPWR VPWR _10801_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12363_ _12363_/A VGND VGND VPWR VPWR _12363_/Y sky130_fd_sc_hd__inv_2
X_15151_ _15134_/A _15134_/B _15134_/Y _15150_/X VGND VGND VPWR VPWR _15151_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14102_ _14098_/Y _14100_/Y _14101_/Y VGND VGND VPWR VPWR _14106_/B sky130_fd_sc_hd__o21ai_1
X_12294_ _13890_/A _12294_/B VGND VGND VPWR VPWR _12294_/X sky130_fd_sc_hd__or2_1
X_15082_ _15082_/A _15028_/X VGND VGND VPWR VPWR _15082_/X sky130_fd_sc_hd__or2b_1
X_11314_ _12268_/A _11314_/B VGND VGND VPWR VPWR _11314_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14033_ _14036_/A VGND VGND VPWR VPWR _15464_/A sky130_fd_sc_hd__buf_1
X_11245_ _12232_/A _13936_/B VGND VGND VPWR VPWR _11245_/X sky130_fd_sc_hd__or2_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11176_ _13894_/A _11176_/B VGND VGND VPWR VPWR _11176_/X sky130_fd_sc_hd__or2_1
XFILLER_79_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15984_ _15984_/A _15984_/B VGND VGND VPWR VPWR _15984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10127_ _10127_/A _10127_/B VGND VGND VPWR VPWR _10128_/B sky130_fd_sc_hd__or2_1
X_14935_ _14835_/X _14849_/A _14848_/X VGND VGND VPWR VPWR _14935_/X sky130_fd_sc_hd__o21a_1
X_10058_ _10019_/X _10057_/Y _10019_/X _10057_/Y VGND VGND VPWR VPWR _10059_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14866_ _14826_/X _14865_/X _14826_/X _14865_/X VGND VGND VPWR VPWR _14926_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14797_ _14730_/X _14796_/X _14730_/X _14796_/X VGND VGND VPWR VPWR _14798_/B sky130_fd_sc_hd__a2bb2o_1
X_13817_ _13764_/X _13816_/X _13764_/X _13816_/X VGND VGND VPWR VPWR _13848_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13748_ _14501_/A _13687_/B _13687_/Y VGND VGND VPWR VPWR _13748_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16467_ _08229_/A _16467_/D VGND VGND VPWR VPWR _16467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13679_ _13618_/X _13678_/X _13618_/X _13678_/X VGND VGND VPWR VPWR _13687_/B sky130_fd_sc_hd__a2bb2o_1
X_16398_ _16407_/B VGND VGND VPWR VPWR _16398_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15418_ _15418_/A _15418_/B VGND VGND VPWR VPWR _15418_/X sky130_fd_sc_hd__or2_1
XFILLER_117_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15349_ _15349_/A _15349_/B VGND VGND VPWR VPWR _15349_/X sky130_fd_sc_hd__or2_1
XFILLER_8_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09910_ _09908_/A _09908_/B _09909_/Y VGND VGND VPWR VPWR _09910_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09841_ _09838_/A _09838_/B _09839_/Y _10500_/A VGND VGND VPWR VPWR _09843_/B sky130_fd_sc_hd__o22a_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09773_/A _09773_/B VGND VGND VPWR VPWR _09772_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08723_ _08843_/A _09459_/B _08719_/Y _08722_/X VGND VGND VPWR VPWR _08723_/X sky130_fd_sc_hd__o22a_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08654_ _08843_/A _09006_/A VGND VGND VPWR VPWR _09799_/A sky130_fd_sc_hd__or2_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08585_ _09467_/B _10115_/B VGND VGND VPWR VPWR _08586_/A sky130_fd_sc_hd__or2_1
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09206_ _13369_/A VGND VGND VPWR VPWR _14012_/A sky130_fd_sc_hd__inv_2
X_09137_ _09133_/Y _09135_/Y _09136_/Y VGND VGND VPWR VPWR _09141_/B sky130_fd_sc_hd__o21ai_1
X_09068_ _10102_/A _09627_/A VGND VGND VPWR VPWR _09069_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11030_ _12846_/A VGND VGND VPWR VPWR _15072_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12981_ _14481_/A _13022_/B VGND VGND VPWR VPWR _13070_/A sky130_fd_sc_hd__and2_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14720_ _11065_/B _14719_/X _11065_/B _14719_/X VGND VGND VPWR VPWR _14722_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11932_ _11912_/X _11931_/X _11912_/X _11931_/X VGND VGND VPWR VPWR _11981_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14651_ _14634_/Y _14649_/X _14650_/Y VGND VGND VPWR VPWR _14651_/X sky130_fd_sc_hd__o21a_1
X_11863_ _12773_/A _11914_/A _11862_/Y VGND VGND VPWR VPWR _11863_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13602_ _13621_/A _13622_/B VGND VGND VPWR VPWR _13602_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10814_ _10078_/X _10813_/X _10078_/X _10813_/X VGND VGND VPWR VPWR _10815_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16321_ _16308_/Y _16319_/X _16320_/Y VGND VGND VPWR VPWR _16321_/X sky130_fd_sc_hd__o21a_1
X_14582_ _14582_/A _14582_/B VGND VGND VPWR VPWR _14582_/Y sky130_fd_sc_hd__nand2_1
X_11794_ _14429_/A _11787_/B _11787_/Y _11793_/X VGND VGND VPWR VPWR _11794_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10745_ _12994_/A _10632_/B _10632_/Y VGND VGND VPWR VPWR _10745_/Y sky130_fd_sc_hd__o21ai_1
X_13533_ _15030_/A _13528_/B _13528_/Y _13532_/X VGND VGND VPWR VPWR _13533_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16252_ _16231_/Y _16250_/X _16251_/Y VGND VGND VPWR VPWR _16252_/X sky130_fd_sc_hd__o21a_1
X_13464_ _15422_/A _12788_/B _12788_/Y _12861_/X VGND VGND VPWR VPWR _13464_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10676_ _10076_/X _10675_/X _10076_/X _10675_/X VGND VGND VPWR VPWR _10677_/B sky130_fd_sc_hd__a2bb2o_1
X_16183_ _15810_/X _16182_/X _15810_/X _16182_/X VGND VGND VPWR VPWR _16184_/B sky130_fd_sc_hd__a2bb2o_1
X_13395_ _14103_/A VGND VGND VPWR VPWR _14106_/A sky130_fd_sc_hd__buf_1
X_15203_ _15137_/A _15137_/B _15137_/Y VGND VGND VPWR VPWR _15203_/Y sky130_fd_sc_hd__o21ai_1
X_12415_ _12679_/A _12426_/B _15560_/A VGND VGND VPWR VPWR _12419_/A sky130_fd_sc_hd__o21ai_2
X_12346_ _12349_/A _12349_/B VGND VGND VPWR VPWR _12346_/Y sky130_fd_sc_hd__nor2_1
X_15134_ _15134_/A _15134_/B VGND VGND VPWR VPWR _15134_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15065_ _15039_/X _15064_/X _15039_/X _15064_/X VGND VGND VPWR VPWR _15066_/B sky130_fd_sc_hd__a2bb2o_1
X_12277_ _12783_/A _12370_/A _12276_/Y VGND VGND VPWR VPWR _12277_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_122_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14016_ _15412_/A _13954_/B _13954_/Y VGND VGND VPWR VPWR _14016_/Y sky130_fd_sc_hd__o21ai_1
X_11228_ _11228_/A _11081_/X VGND VGND VPWR VPWR _11228_/X sky130_fd_sc_hd__or2b_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ _11139_/X _11158_/X _11139_/X _11158_/X VGND VGND VPWR VPWR _11304_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15967_ _15906_/A _15906_/B _15906_/Y VGND VGND VPWR VPWR _15967_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15898_ _15898_/A _15898_/B VGND VGND VPWR VPWR _15898_/Y sky130_fd_sc_hd__nand2_1
X_14918_ _15542_/A _14918_/B VGND VGND VPWR VPWR _14918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14849_ _14849_/A _14848_/X VGND VGND VPWR VPWR _14849_/X sky130_fd_sc_hd__or2b_1
XFILLER_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ _08263_/A input14/X _08342_/B _08418_/A VGND VGND VPWR VPWR _08424_/A sky130_fd_sc_hd__o22a_1
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09824_ _09819_/A _09819_/B _09820_/B VGND VGND VPWR VPWR _09843_/A sky130_fd_sc_hd__a21bo_1
XFILLER_100_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09742_/A _09742_/B _09745_/A VGND VGND VPWR VPWR _10085_/A sky130_fd_sc_hd__a21bo_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08706_ _09341_/A _08706_/B VGND VGND VPWR VPWR _08749_/A sky130_fd_sc_hd__or2_2
X_09686_ _09686_/A _09686_/B VGND VGND VPWR VPWR _09689_/A sky130_fd_sc_hd__or2_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08637_ _08637_/A VGND VGND VPWR VPWR _08637_/Y sky130_fd_sc_hd__inv_2
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08567_/X _08433_/X _08567_/X _08433_/X VGND VGND VPWR VPWR _08571_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08499_ _08650_/A VGND VGND VPWR VPWR _08589_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10530_ _10497_/Y _10528_/X _10529_/Y VGND VGND VPWR VPWR _10530_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10461_ _10461_/A VGND VGND VPWR VPWR _10461_/Y sky130_fd_sc_hd__inv_2
X_12200_ _13894_/A _12200_/B VGND VGND VPWR VPWR _12200_/X sky130_fd_sc_hd__or2_1
X_13180_ _14568_/A _13101_/B _13101_/Y VGND VGND VPWR VPWR _13180_/Y sky130_fd_sc_hd__o21ai_1
X_10392_ _11770_/A _10392_/B VGND VGND VPWR VPWR _10392_/X sky130_fd_sc_hd__and2_1
XFILLER_108_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12131_ _12137_/A _12137_/B VGND VGND VPWR VPWR _12228_/A sky130_fd_sc_hd__and2_1
XFILLER_123_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12062_ _12018_/Y _12060_/X _12061_/Y VGND VGND VPWR VPWR _12062_/X sky130_fd_sc_hd__o21a_1
X_11013_ _13902_/A _11091_/B VGND VGND VPWR VPWR _11195_/A sky130_fd_sc_hd__and2_1
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15821_ _16123_/A _15821_/B VGND VGND VPWR VPWR _16142_/B sky130_fd_sc_hd__or2_1
XFILLER_77_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15752_ _15752_/A _15752_/B VGND VGND VPWR VPWR _16106_/A sky130_fd_sc_hd__nor2_1
XFILLER_92_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12964_ _12941_/X _12963_/Y _12941_/X _12963_/Y VGND VGND VPWR VPWR _13030_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14703_ _15339_/A _14654_/B _14654_/Y VGND VGND VPWR VPWR _14703_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11915_ _11913_/A _11913_/B _11913_/X _11914_/Y VGND VGND VPWR VPWR _11985_/B sky130_fd_sc_hd__a22o_1
XFILLER_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15683_ _15683_/A _15683_/B VGND VGND VPWR VPWR _15683_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12895_ _14467_/A _12932_/B VGND VGND VPWR VPWR _12895_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _15335_/A _14650_/B VGND VGND VPWR VPWR _14634_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11846_ _13556_/A _11845_/B _11845_/X _11797_/X VGND VGND VPWR VPWR _11846_/X sky130_fd_sc_hd__o22a_1
XFILLER_54_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _14565_/A _14510_/X VGND VGND VPWR VPWR _14565_/X sky130_fd_sc_hd__or2b_1
X_11777_ _12765_/A _11777_/B VGND VGND VPWR VPWR _11777_/Y sky130_fd_sc_hd__nor2_1
X_16304_ _16254_/X _16303_/Y _16254_/X _16303_/Y VGND VGND VPWR VPWR _16322_/B sky130_fd_sc_hd__o2bb2a_1
X_10728_ _10637_/A _10727_/Y _10637_/A _10727_/Y VGND VGND VPWR VPWR _10729_/B sky130_fd_sc_hd__a2bb2o_1
X_13516_ _13516_/A _13516_/B VGND VGND VPWR VPWR _13516_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16235_ _16233_/A _16234_/A _16233_/Y _16234_/Y _16243_/A VGND VGND VPWR VPWR _16249_/A
+ sky130_fd_sc_hd__a221o_1
X_14496_ _15205_/A _14514_/B VGND VGND VPWR VPWR _14557_/A sky130_fd_sc_hd__and2_1
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13447_ _13381_/Y _13445_/X _13446_/Y VGND VGND VPWR VPWR _13447_/X sky130_fd_sc_hd__o21a_1
X_10659_ _09269_/A _09269_/B _09269_/X VGND VGND VPWR VPWR _10660_/B sky130_fd_sc_hd__a21boi_1
X_16166_ _16114_/A _15815_/B _15815_/Y VGND VGND VPWR VPWR _16166_/X sky130_fd_sc_hd__o21a_1
X_13378_ _14144_/A _13448_/B VGND VGND VPWR VPWR _13378_/Y sky130_fd_sc_hd__nor2_1
X_16097_ _16034_/A _16034_/B _16034_/Y VGND VGND VPWR VPWR _16097_/Y sky130_fd_sc_hd__o21ai_1
X_12329_ _12329_/A _12329_/B VGND VGND VPWR VPWR _12329_/X sky130_fd_sc_hd__or2_1
X_15117_ _15060_/A _15060_/B _15060_/Y VGND VGND VPWR VPWR _15117_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15048_ _12180_/A _15006_/X _12179_/X VGND VGND VPWR VPWR _15048_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09540_ _09540_/A _09540_/B VGND VGND VPWR VPWR _09540_/X sky130_fd_sc_hd__or2_1
XFILLER_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09471_ _09452_/Y _09469_/X _09470_/X VGND VGND VPWR VPWR _09471_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08422_ _08715_/A VGND VGND VPWR VPWR _09250_/A sky130_fd_sc_hd__buf_1
XFILLER_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08353_ _08353_/A _08353_/B VGND VGND VPWR VPWR _08354_/A sky130_fd_sc_hd__or2_1
XFILLER_20_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08284_ input26/X _08357_/B _08387_/A _08389_/A VGND VGND VPWR VPWR _08384_/A sky130_fd_sc_hd__o22a_1
XFILLER_109_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09807_ _08852_/A _08721_/B _09817_/A VGND VGND VPWR VPWR _09808_/A sky130_fd_sc_hd__o21ai_1
XFILLER_86_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09738_ _08546_/A _09740_/B _08546_/A _09740_/B VGND VGND VPWR VPWR _09739_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09562_/Y _09668_/Y _09562_/Y _09668_/Y VGND VGND VPWR VPWR _09669_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_82_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _15556_/A _11641_/B _11641_/X _11644_/Y VGND VGND VPWR VPWR _11700_/X sky130_fd_sc_hd__a22o_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12680_ _12425_/A _12679_/B _12679_/Y VGND VGND VPWR VPWR _12680_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _12440_/A _11631_/B VGND VGND VPWR VPWR _11631_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14350_ _14253_/A _14349_/Y _14253_/A _14349_/Y VGND VGND VPWR VPWR _14380_/A sky130_fd_sc_hd__a2bb2o_1
X_11562_ _14066_/A _11561_/B _11561_/Y VGND VGND VPWR VPWR _11562_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13301_ _13225_/Y _13299_/Y _13300_/Y VGND VGND VPWR VPWR _13302_/A sky130_fd_sc_hd__o21ai_1
X_10513_ _10431_/X _10512_/X _10431_/X _10512_/X VGND VGND VPWR VPWR _10525_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14281_ _14134_/X _14280_/Y _14134_/X _14280_/Y VGND VGND VPWR VPWR _14282_/B sky130_fd_sc_hd__a2bb2oi_1
X_11493_ _11491_/Y _11492_/Y _11341_/Y VGND VGND VPWR VPWR _11493_/X sky130_fd_sc_hd__o21a_1
X_16020_ _16020_/A _15950_/X VGND VGND VPWR VPWR _16020_/X sky130_fd_sc_hd__or2b_1
X_13232_ _14529_/A VGND VGND VPWR VPWR _14737_/A sky130_fd_sc_hd__buf_1
X_10444_ _09978_/A _09978_/B _09978_/Y VGND VGND VPWR VPWR _10445_/A sky130_fd_sc_hd__o21ai_1
XFILLER_123_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13163_ _15255_/A _13111_/B _13111_/Y VGND VGND VPWR VPWR _13163_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10375_ _10251_/A _10170_/B _10170_/Y VGND VGND VPWR VPWR _10376_/A sky130_fd_sc_hd__a21oi_1
XFILLER_124_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12114_ _13194_/A _12059_/B _12059_/Y VGND VGND VPWR VPWR _12114_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13094_ _13009_/X _13093_/Y _13009_/X _13093_/Y VGND VGND VPWR VPWR _13103_/B sky130_fd_sc_hd__a2bb2o_1
X_12045_ _11062_/A _12044_/X _11062_/A _12044_/X VGND VGND VPWR VPWR _12047_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15804_ _15672_/X _15803_/Y _15672_/X _15803_/Y VGND VGND VPWR VPWR _16207_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13996_ _13963_/X _13994_/Y _13995_/Y VGND VGND VPWR VPWR _13996_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15735_ _15681_/A _15681_/B _15681_/Y VGND VGND VPWR VPWR _15735_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12947_ _14944_/A _12947_/B VGND VGND VPWR VPWR _12947_/Y sky130_fd_sc_hd__nand2_1
X_15666_ _15774_/A _16028_/A _15775_/B _15665_/X VGND VGND VPWR VPWR _15666_/X sky130_fd_sc_hd__a31o_1
XFILLER_73_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12878_ _12853_/X _12877_/Y _12853_/X _12877_/Y VGND VGND VPWR VPWR _12940_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14617_ _14585_/X _14616_/Y _14585_/X _14616_/Y VGND VGND VPWR VPWR _14658_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11829_ _11793_/X _11828_/X _11793_/X _11828_/X VGND VGND VPWR VPWR _11835_/B sky130_fd_sc_hd__a2bb2o_1
X_15597_ _15597_/A _14392_/X VGND VGND VPWR VPWR _15597_/X sky130_fd_sc_hd__or2b_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14548_ _15255_/A VGND VGND VPWR VPWR _14582_/A sky130_fd_sc_hd__buf_1
X_14479_ _14470_/X _14478_/X _14470_/X _14478_/X VGND VGND VPWR VPWR _14522_/B sky130_fd_sc_hd__a2bb2o_1
X_16218_ _16218_/A VGND VGND VPWR VPWR _16218_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16149_ _16147_/A _16148_/A _16147_/Y _16148_/Y _16388_/A VGND VGND VPWR VPWR _16270_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08971_ _08912_/X _08969_/X _11389_/B VGND VGND VPWR VPWR _08971_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09523_ _09521_/Y _09522_/X _09521_/Y _09522_/X VGND VGND VPWR VPWR _09523_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09454_ _09492_/A _09454_/B VGND VGND VPWR VPWR _09454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08405_ _08653_/A VGND VGND VPWR VPWR _08944_/A sky130_fd_sc_hd__inv_2
X_09385_ _09432_/B _09383_/B _09383_/X _11096_/A VGND VGND VPWR VPWR _11269_/A sky130_fd_sc_hd__a22o_1
XFILLER_51_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08336_ _08336_/A input31/X VGND VGND VPWR VPWR _08337_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08267_ input12/X VGND VGND VPWR VPWR _08352_/B sky130_fd_sc_hd__inv_2
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10160_ _10114_/A _10114_/B _10115_/A VGND VGND VPWR VPWR _10163_/A sky130_fd_sc_hd__a21bo_1
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10091_ _09194_/Y _10090_/X _09194_/Y _10090_/X VGND VGND VPWR VPWR _10091_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13850_ _14619_/A _13850_/B VGND VGND VPWR VPWR _13850_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13781_ _13789_/A VGND VGND VPWR VPWR _15113_/A sky130_fd_sc_hd__buf_1
X_10993_ _13706_/A _11122_/B _10992_/Y VGND VGND VPWR VPWR _10993_/Y sky130_fd_sc_hd__o21ai_1
X_12801_ _12854_/A _12854_/B VGND VGND VPWR VPWR _12801_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15520_ _15639_/A _15640_/A _15519_/X VGND VGND VPWR VPWR _15524_/B sky130_fd_sc_hd__o21ai_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12781_/A _12781_/B VGND VGND VPWR VPWR _12732_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15451_ _15409_/X _15450_/X _15409_/X _15450_/X VGND VGND VPWR VPWR _15452_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14402_ _15687_/A _14400_/Y _14401_/X VGND VGND VPWR VPWR _14402_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12663_ _10554_/Y _12662_/Y _10465_/Y VGND VGND VPWR VPWR _12664_/A sky130_fd_sc_hd__o21ai_1
X_12594_ _12594_/A VGND VGND VPWR VPWR _12594_/Y sky130_fd_sc_hd__inv_2
X_15382_ _15336_/X _15381_/X _15336_/X _15381_/X VGND VGND VPWR VPWR _15404_/B sky130_fd_sc_hd__a2bb2o_1
X_11614_ _11611_/X _11689_/A _11611_/A _11689_/A VGND VGND VPWR VPWR _11615_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_128_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14333_ _14106_/A _13431_/B _13431_/Y VGND VGND VPWR VPWR _14333_/X sky130_fd_sc_hd__o21a_1
X_11545_ _11499_/X _11544_/Y _11499_/X _11544_/Y VGND VGND VPWR VPWR _11643_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14264_ _14210_/Y _14262_/Y _14263_/Y VGND VGND VPWR VPWR _14265_/A sky130_fd_sc_hd__o21ai_2
X_11476_ _12440_/A VGND VGND VPWR VPWR _13872_/A sky130_fd_sc_hd__buf_1
XFILLER_51_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16003_ _15961_/X _16002_/X _15961_/X _16002_/X VGND VGND VPWR VPWR _16044_/B sky130_fd_sc_hd__a2bb2o_1
X_13215_ _14858_/A _13306_/B VGND VGND VPWR VPWR _13215_/Y sky130_fd_sc_hd__nor2_1
X_10427_ _12232_/A _11792_/B VGND VGND VPWR VPWR _10622_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14195_ _14207_/A _14195_/B VGND VGND VPWR VPWR _15863_/A sky130_fd_sc_hd__or2_1
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13146_ _13122_/X _13145_/Y _13122_/X _13145_/Y VGND VGND VPWR VPWR _13204_/B sky130_fd_sc_hd__a2bb2o_1
X_10358_ _15028_/A _10338_/B _10338_/X _10357_/X VGND VGND VPWR VPWR _10358_/X sky130_fd_sc_hd__o22a_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13077_ _15255_/A _13111_/B VGND VGND VPWR VPWR _13077_/Y sky130_fd_sc_hd__nor2_1
X_10289_ _10289_/A _10352_/A VGND VGND VPWR VPWR _10289_/X sky130_fd_sc_hd__or2_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12028_ _13078_/A _11970_/B _11970_/Y VGND VGND VPWR VPWR _12028_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13979_ _13979_/A _13979_/B VGND VGND VPWR VPWR _13979_/X sky130_fd_sc_hd__or2_1
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15718_ _16121_/A _15819_/B VGND VGND VPWR VPWR _15718_/X sky130_fd_sc_hd__and2_1
XFILLER_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15649_ _15512_/A _15512_/B _15512_/X VGND VGND VPWR VPWR _15650_/A sky130_fd_sc_hd__o21ba_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09170_ _09750_/A VGND VGND VPWR VPWR _09429_/A sky130_fd_sc_hd__buf_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08954_ _10018_/A _10124_/A _08836_/Y VGND VGND VPWR VPWR _08954_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08885_ _08980_/A _08980_/B VGND VGND VPWR VPWR _08885_/X sky130_fd_sc_hd__and2_1
XFILLER_29_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09506_ _08922_/A _09503_/Y _09503_/A _09505_/Y VGND VGND VPWR VPWR _09506_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09437_ _09323_/A _09435_/Y _09436_/Y VGND VGND VPWR VPWR _11106_/A sky130_fd_sc_hd__o21ai_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ _09368_/A VGND VGND VPWR VPWR _09430_/B sky130_fd_sc_hd__inv_2
X_09299_ _09299_/A VGND VGND VPWR VPWR _09299_/Y sky130_fd_sc_hd__inv_2
X_08319_ _08319_/A VGND VGND VPWR VPWR _08319_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11330_ _11329_/A _11329_/B _11329_/Y _10982_/X VGND VGND VPWR VPWR _12373_/A sky130_fd_sc_hd__o211a_1
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11261_ _15443_/A _11179_/B _11179_/Y _11260_/X VGND VGND VPWR VPWR _11261_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11192_ _13365_/A VGND VGND VPWR VPWR _14018_/A sky130_fd_sc_hd__inv_2
X_13000_ _13677_/A _13010_/B VGND VGND VPWR VPWR _13000_/Y sky130_fd_sc_hd__nor2_1
X_10212_ _10282_/A _11721_/A _10281_/A VGND VGND VPWR VPWR _10212_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10143_ _10143_/A _10143_/B VGND VGND VPWR VPWR _10143_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14951_ _14976_/A _14976_/B VGND VGND VPWR VPWR _14951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10074_ _10023_/X _10073_/Y _10023_/X _10073_/Y VGND VGND VPWR VPWR _10075_/B sky130_fd_sc_hd__a2bb2o_1
X_14882_ _14822_/X _14881_/X _14822_/X _14881_/X VGND VGND VPWR VPWR _14918_/B sky130_fd_sc_hd__a2bb2o_1
X_13902_ _13902_/A VGND VGND VPWR VPWR _15412_/A sky130_fd_sc_hd__buf_1
XFILLER_75_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13833_ _13833_/A VGND VGND VPWR VPWR _13838_/A sky130_fd_sc_hd__inv_2
XFILLER_75_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15503_ _15544_/A _15544_/B VGND VGND VPWR VPWR _15503_/X sky130_fd_sc_hd__and2_1
X_13764_ _13819_/A _13762_/X _13763_/X VGND VGND VPWR VPWR _13764_/X sky130_fd_sc_hd__o21a_1
X_10976_ _12174_/A _11140_/B VGND VGND VPWR VPWR _10976_/Y sky130_fd_sc_hd__nand2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13695_ _13695_/A _13695_/B VGND VGND VPWR VPWR _13695_/X sky130_fd_sc_hd__or2_1
X_12715_ _12692_/A _12692_/B _12692_/Y _12714_/X VGND VGND VPWR VPWR _12715_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12646_ _14984_/A _12494_/B _12494_/Y VGND VGND VPWR VPWR _12646_/X sky130_fd_sc_hd__o21a_1
X_15434_ _15563_/A _15563_/B _15433_/Y VGND VGND VPWR VPWR _15434_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15365_ _15416_/A _15416_/B VGND VGND VPWR VPWR _15441_/A sky130_fd_sc_hd__and2_1
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14316_ _15860_/A _14272_/B _14272_/Y VGND VGND VPWR VPWR _14316_/Y sky130_fd_sc_hd__o21ai_1
X_12577_ _14910_/A _11434_/B _11434_/Y VGND VGND VPWR VPWR _12578_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15296_ _15351_/A _15351_/B VGND VGND VPWR VPWR _15360_/A sky130_fd_sc_hd__and2_1
X_11528_ _11528_/A _11528_/B VGND VGND VPWR VPWR _11528_/X sky130_fd_sc_hd__or2_1
XFILLER_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14247_ _11705_/A _14362_/B _12500_/A _15778_/A VGND VGND VPWR VPWR _15838_/A sky130_fd_sc_hd__o22a_1
X_11459_ _14138_/A _11356_/B _11356_/Y _12506_/A VGND VGND VPWR VPWR _11566_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14178_ _14178_/A _12635_/X VGND VGND VPWR VPWR _14178_/X sky130_fd_sc_hd__or2b_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13129_ _12952_/A _13035_/X _12951_/X VGND VGND VPWR VPWR _13129_/X sky130_fd_sc_hd__o21a_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08670_ _08670_/A VGND VGND VPWR VPWR _08929_/A sky130_fd_sc_hd__inv_2
XFILLER_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09222_ _09802_/A VGND VGND VPWR VPWR _09693_/A sky130_fd_sc_hd__inv_2
XFILLER_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09153_ _08762_/A _09147_/X _09147_/X _08535_/Y VGND VGND VPWR VPWR _09154_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09084_ _09766_/A VGND VGND VPWR VPWR _09426_/A sky130_fd_sc_hd__buf_1
XFILLER_116_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09986_ _09986_/A _09987_/B VGND VGND VPWR VPWR _09986_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08937_ _09041_/A _08937_/B VGND VGND VPWR VPWR _08937_/X sky130_fd_sc_hd__or2_1
X_08868_ _09482_/A _08760_/Y _08762_/Y _08867_/X VGND VGND VPWR VPWR _08868_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08799_ _08798_/X _08731_/Y _08798_/A _08731_/Y VGND VGND VPWR VPWR _08801_/A sky130_fd_sc_hd__a2bb2o_1
X_10830_ _10962_/A _12690_/A _10829_/Y VGND VGND VPWR VPWR _10830_/X sky130_fd_sc_hd__a21o_1
X_10761_ _10761_/A _12605_/A VGND VGND VPWR VPWR _13754_/A sky130_fd_sc_hd__or2_1
XFILLER_53_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12500_ _12500_/A VGND VGND VPWR VPWR _12501_/A sky130_fd_sc_hd__clkbuf_2
X_13480_ _10421_/B _13479_/Y _11713_/A _10286_/B VGND VGND VPWR VPWR _13481_/A sky130_fd_sc_hd__o22a_1
X_10692_ _10809_/A _12692_/A _10691_/Y VGND VGND VPWR VPWR _10692_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12431_ _13458_/A _12421_/Y _12429_/A _12428_/X _12430_/X VGND VGND VPWR VPWR _12431_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_40_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12362_ _12362_/A _12362_/B VGND VGND VPWR VPWR _12362_/Y sky130_fd_sc_hd__nor2_1
X_15150_ _15137_/A _15137_/B _15137_/Y _15149_/X VGND VGND VPWR VPWR _15150_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14101_ _14101_/A _14101_/B VGND VGND VPWR VPWR _14101_/Y sky130_fd_sc_hd__nand2_1
X_12293_ _13890_/A _12294_/B VGND VGND VPWR VPWR _12295_/A sky130_fd_sc_hd__and2_1
X_15081_ _15081_/A _15081_/B VGND VGND VPWR VPWR _15081_/Y sky130_fd_sc_hd__nand2_1
X_11313_ _11309_/Y _12686_/A _11139_/X _11312_/Y VGND VGND VPWR VPWR _11313_/X sky130_fd_sc_hd__o22a_1
X_14032_ _14032_/A _14032_/B VGND VGND VPWR VPWR _14032_/X sky130_fd_sc_hd__and2_1
X_11244_ _11244_/A VGND VGND VPWR VPWR _13936_/B sky130_fd_sc_hd__buf_1
XFILLER_4_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11175_ _13894_/A _11176_/B VGND VGND VPWR VPWR _11177_/A sky130_fd_sc_hd__and2_1
X_15983_ _15973_/X _15988_/A _15982_/X VGND VGND VPWR VPWR _15983_/Y sky130_fd_sc_hd__o21ai_1
X_10126_ _10126_/A _10126_/B VGND VGND VPWR VPWR _10127_/B sky130_fd_sc_hd__or2_1
XFILLER_94_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14934_ _14934_/A VGND VGND VPWR VPWR _14971_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10057_ _08843_/A _09070_/A _08944_/X VGND VGND VPWR VPWR _10057_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14865_ _14774_/A _14774_/B _14774_/A _14774_/B VGND VGND VPWR VPWR _14865_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14796_ _14796_/A _14731_/X VGND VGND VPWR VPWR _14796_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13816_ _13816_/A _13765_/X VGND VGND VPWR VPWR _13816_/X sky130_fd_sc_hd__or2b_1
X_13747_ _13747_/A _13759_/B VGND VGND VPWR VPWR _13826_/A sky130_fd_sc_hd__and2_1
X_10959_ _12078_/A VGND VGND VPWR VPWR _13507_/A sky130_fd_sc_hd__buf_1
X_16466_ _16357_/A _16466_/D VGND VGND VPWR VPWR _16466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15417_ _15441_/A _15415_/X _15416_/X VGND VGND VPWR VPWR _15417_/X sky130_fd_sc_hd__o21a_1
X_13678_ _12923_/A _13609_/B _12923_/A _13609_/B VGND VGND VPWR VPWR _13678_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16397_ _16397_/A _16397_/B _16397_/C _16397_/D VGND VGND VPWR VPWR _16407_/B sky130_fd_sc_hd__or4_1
XFILLER_129_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12629_ _12629_/A _12629_/B VGND VGND VPWR VPWR _12629_/X sky130_fd_sc_hd__or2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15348_ _15366_/A _15346_/X _15347_/X VGND VGND VPWR VPWR _15348_/X sky130_fd_sc_hd__o21a_1
X_15279_ _14586_/A _15249_/B _15249_/Y _15278_/X VGND VGND VPWR VPWR _15279_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _09687_/A _09834_/Y _09801_/B VGND VGND VPWR VPWR _10500_/A sky130_fd_sc_hd__o21ai_2
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09700_/A _09770_/Y _09725_/Y VGND VGND VPWR VPWR _09773_/B sky130_fd_sc_hd__o21ai_2
X_08722_ _08852_/A _09540_/A _09235_/A _09041_/A VGND VGND VPWR VPWR _08722_/X sky130_fd_sc_hd__o22a_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08653_ _08653_/A VGND VGND VPWR VPWR _08843_/A sky130_fd_sc_hd__buf_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08584_ _08584_/A VGND VGND VPWR VPWR _10115_/B sky130_fd_sc_hd__inv_2
XFILLER_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09205_ _09040_/Y _09145_/A _09040_/A _09145_/Y _09204_/X VGND VGND VPWR VPWR _13369_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_10_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09136_ _09426_/A _09136_/B VGND VGND VPWR VPWR _09136_/Y sky130_fd_sc_hd__nand2_1
X_09067_ _08930_/A _09829_/A _08922_/A VGND VGND VPWR VPWR _09627_/A sky130_fd_sc_hd__o21ai_2
XFILLER_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09969_ _10077_/A VGND VGND VPWR VPWR _09969_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12980_ _12933_/X _12979_/Y _12933_/X _12979_/Y VGND VGND VPWR VPWR _13022_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11931_ _11014_/A _11983_/B _11014_/A _11983_/B VGND VGND VPWR VPWR _11931_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14650_ _15335_/A _14650_/B VGND VGND VPWR VPWR _14650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11862_ _12773_/A _11914_/A VGND VGND VPWR VPWR _11862_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14581_ _14555_/Y _14579_/X _14580_/Y VGND VGND VPWR VPWR _14581_/X sky130_fd_sc_hd__o21a_1
X_13601_ _13576_/X _13600_/Y _13576_/X _13600_/Y VGND VGND VPWR VPWR _13622_/B sky130_fd_sc_hd__a2bb2o_1
X_10813_ _10049_/X _10813_/B VGND VGND VPWR VPWR _10813_/X sky130_fd_sc_hd__and2b_1
X_16320_ _16320_/A _16320_/B VGND VGND VPWR VPWR _16320_/Y sky130_fd_sc_hd__nand2_1
X_11793_ _12826_/A _11791_/B _11791_/X _11792_/X VGND VGND VPWR VPWR _11793_/X sky130_fd_sc_hd__o22a_1
X_13532_ _15028_/A _13530_/B _13530_/Y _13531_/X VGND VGND VPWR VPWR _13532_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10744_ _10744_/A VGND VGND VPWR VPWR _12994_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16251_ _16251_/A _16251_/B VGND VGND VPWR VPWR _16251_/Y sky130_fd_sc_hd__nand2_1
X_13463_ _13463_/A VGND VGND VPWR VPWR _15422_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10675_ _10052_/X _10675_/B VGND VGND VPWR VPWR _10675_/X sky130_fd_sc_hd__and2b_1
X_16182_ _16110_/A _15811_/B _15811_/Y VGND VGND VPWR VPWR _16182_/X sky130_fd_sc_hd__o21a_1
X_13394_ _14108_/A VGND VGND VPWR VPWR _14112_/A sky130_fd_sc_hd__buf_1
X_15202_ _15202_/A _15202_/B VGND VGND VPWR VPWR _15202_/Y sky130_fd_sc_hd__nand2_1
X_12414_ _12679_/A _12426_/B VGND VGND VPWR VPWR _15560_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12345_ _12341_/Y _12559_/A _12344_/Y VGND VGND VPWR VPWR _12349_/B sky130_fd_sc_hd__o21ai_1
X_15133_ _15091_/X _15132_/Y _15091_/X _15132_/Y VGND VGND VPWR VPWR _15134_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12276_ _12369_/A _12370_/A VGND VGND VPWR VPWR _12276_/Y sky130_fd_sc_hd__nor2_1
X_15064_ _15064_/A _15040_/X VGND VGND VPWR VPWR _15064_/X sky130_fd_sc_hd__or2b_1
X_11227_ _12224_/A VGND VGND VPWR VPWR _14036_/A sky130_fd_sc_hd__buf_1
X_14015_ _14015_/A _14060_/B VGND VGND VPWR VPWR _14123_/A sky130_fd_sc_hd__and2_1
XFILLER_110_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11158_ _11312_/A _12266_/A _11157_/Y VGND VGND VPWR VPWR _11158_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10109_ _10109_/A VGND VGND VPWR VPWR _10109_/Y sky130_fd_sc_hd__inv_2
X_15966_ _15966_/A _15966_/B VGND VGND VPWR VPWR _15966_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11089_ _13906_/A _11089_/B VGND VGND VPWR VPWR _11089_/X sky130_fd_sc_hd__or2_1
XFILLER_76_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15897_ _15868_/Y _15895_/X _15896_/Y VGND VGND VPWR VPWR _15897_/X sky130_fd_sc_hd__o21a_1
X_14917_ _14886_/Y _14915_/X _14916_/Y VGND VGND VPWR VPWR _14917_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14848_ _15178_/A _14848_/B VGND VGND VPWR VPWR _14848_/X sky130_fd_sc_hd__or2_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14779_ _15446_/A VGND VGND VPWR VPWR _14782_/A sky130_fd_sc_hd__buf_1
XFILLER_90_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16449_ _16412_/Y _16473_/Q _16446_/Y _16428_/Y VGND VGND VPWR VPWR _16449_/X sky130_fd_sc_hd__o211a_1
XFILLER_129_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09823_ _09820_/A _09820_/B _09821_/B VGND VGND VPWR VPWR _09848_/A sky130_fd_sc_hd__a21bo_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _09754_/A VGND VGND VPWR VPWR _09788_/A sky130_fd_sc_hd__inv_2
XFILLER_67_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08705_ _09342_/A VGND VGND VPWR VPWR _08706_/B sky130_fd_sc_hd__inv_2
X_09685_ _08645_/X _09687_/B _08645_/A _09687_/B VGND VGND VPWR VPWR _09686_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08636_ _09462_/B _10111_/B VGND VGND VPWR VPWR _08637_/A sky130_fd_sc_hd__or2_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08567_ _09734_/A _08567_/B VGND VGND VPWR VPWR _08567_/X sky130_fd_sc_hd__or2_1
XFILLER_120_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08498_ _08660_/A VGND VGND VPWR VPWR _08650_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10460_ _10469_/A _10167_/B _10167_/Y VGND VGND VPWR VPWR _10461_/A sky130_fd_sc_hd__a21oi_1
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09119_ _09115_/Y _09117_/Y _09118_/Y VGND VGND VPWR VPWR _09123_/B sky130_fd_sc_hd__o21ai_1
XFILLER_89_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10391_ _10360_/X _10390_/X _10360_/X _10390_/X VGND VGND VPWR VPWR _10392_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12130_ _12048_/X _12129_/Y _12048_/X _12129_/Y VGND VGND VPWR VPWR _12137_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12061_ _12061_/A _12061_/B VGND VGND VPWR VPWR _12061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11012_ _10920_/X _11011_/X _10920_/X _11011_/X VGND VGND VPWR VPWR _11091_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15820_ _15718_/X _15818_/X _16150_/B VGND VGND VPWR VPWR _15820_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15751_ _14913_/X _15750_/X _14913_/X _15750_/X VGND VGND VPWR VPWR _15752_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_73_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12963_ _14677_/A _12942_/B _12942_/Y VGND VGND VPWR VPWR _12963_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15682_ _15599_/Y _15680_/X _15681_/Y VGND VGND VPWR VPWR _15682_/X sky130_fd_sc_hd__o21a_1
X_14702_ _14733_/A _14733_/B VGND VGND VPWR VPWR _14792_/A sky130_fd_sc_hd__and2_1
X_11914_ _11914_/A VGND VGND VPWR VPWR _11914_/Y sky130_fd_sc_hd__inv_2
X_14633_ _14577_/X _14632_/Y _14577_/X _14632_/Y VGND VGND VPWR VPWR _14650_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12894_ _12845_/X _12893_/Y _12845_/X _12893_/Y VGND VGND VPWR VPWR _12932_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _13556_/A _11845_/B VGND VGND VPWR VPWR _11845_/X sky130_fd_sc_hd__and2_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14564_/A VGND VGND VPWR VPWR _15272_/A sky130_fd_sc_hd__buf_1
X_11776_ _11776_/A VGND VGND VPWR VPWR _12765_/A sky130_fd_sc_hd__buf_1
XFILLER_14_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16303_ _16255_/A _16322_/A _16255_/Y VGND VGND VPWR VPWR _16303_/Y sky130_fd_sc_hd__o21ai_1
X_14495_ _14462_/X _14494_/Y _14462_/X _14494_/Y VGND VGND VPWR VPWR _14514_/B sky130_fd_sc_hd__a2bb2o_1
X_10727_ _13693_/A _10638_/B _10638_/Y VGND VGND VPWR VPWR _10727_/Y sky130_fd_sc_hd__o21ai_1
X_13515_ _10573_/X _13486_/X _10573_/X _13486_/X VGND VGND VPWR VPWR _13516_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16234_ _16234_/A VGND VGND VPWR VPWR _16234_/Y sky130_fd_sc_hd__inv_2
X_13446_ _13446_/A _13446_/B VGND VGND VPWR VPWR _13446_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10658_ _10543_/X _10657_/B _10657_/X _10539_/X VGND VGND VPWR VPWR _10658_/X sky130_fd_sc_hd__o22a_1
XFILLER_127_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16165_ _16189_/A _16165_/B VGND VGND VPWR VPWR _16266_/A sky130_fd_sc_hd__or2_1
X_13377_ _13372_/X _13376_/X _13372_/X _13376_/X VGND VGND VPWR VPWR _13448_/B sky130_fd_sc_hd__a2bb2o_1
X_10589_ _09720_/A _09720_/B _09720_/Y VGND VGND VPWR VPWR _10590_/A sky130_fd_sc_hd__o21ai_1
X_16096_ _16099_/A _16099_/B VGND VGND VPWR VPWR _16096_/Y sky130_fd_sc_hd__nor2_1
X_12328_ _12238_/X _12327_/Y _12238_/X _12327_/Y VGND VGND VPWR VPWR _12589_/A sky130_fd_sc_hd__a2bb2o_1
X_15116_ _15116_/A _15116_/B VGND VGND VPWR VPWR _15116_/Y sky130_fd_sc_hd__nand2_1
X_12259_ _12259_/A _12259_/B VGND VGND VPWR VPWR _12259_/X sky130_fd_sc_hd__and2_1
X_15047_ _15055_/A _15045_/X _15046_/X VGND VGND VPWR VPWR _15047_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15949_ _16023_/A _15947_/Y _15948_/X VGND VGND VPWR VPWR _15949_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09470_ _09470_/A _09470_/B VGND VGND VPWR VPWR _09470_/X sky130_fd_sc_hd__or2_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08421_ _09217_/A VGND VGND VPWR VPWR _08715_/A sky130_fd_sc_hd__inv_2
XFILLER_17_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08352_ input28/X _08352_/B VGND VGND VPWR VPWR _08353_/B sky130_fd_sc_hd__nor2_1
X_08283_ _08276_/Y input25/X _08279_/Y _08399_/B VGND VGND VPWR VPWR _08389_/A sky130_fd_sc_hd__o22a_1
XFILLER_20_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09806_ _09855_/B VGND VGND VPWR VPWR _09806_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09737_ _09737_/A _09737_/B VGND VGND VPWR VPWR _09740_/B sky130_fd_sc_hd__or2_1
XFILLER_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09668_ _09569_/A _09569_/B _09569_/Y _09667_/Y VGND VGND VPWR VPWR _09668_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09599_ _09511_/X _09598_/X _09511_/X _09598_/X VGND VGND VPWR VPWR _09983_/A sky130_fd_sc_hd__a2bb2o_1
X_08619_ _08618_/X _08413_/Y _08618_/X _08413_/Y VGND VGND VPWR VPWR _08622_/A sky130_fd_sc_hd__o2bb2a_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11630_ _13133_/A _11629_/B _11629_/Y VGND VGND VPWR VPWR _11630_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11561_ _14066_/A _11561_/B VGND VGND VPWR VPWR _11561_/Y sky130_fd_sc_hd__nand2_1
X_13300_ _14741_/A _13300_/B VGND VGND VPWR VPWR _13300_/Y sky130_fd_sc_hd__nand2_1
X_10512_ _10512_/A _10432_/X VGND VGND VPWR VPWR _10512_/X sky130_fd_sc_hd__or2b_1
X_14280_ _13446_/A _14139_/A _14137_/Y VGND VGND VPWR VPWR _14280_/Y sky130_fd_sc_hd__a21oi_1
X_11492_ _11492_/A VGND VGND VPWR VPWR _11492_/Y sky130_fd_sc_hd__inv_2
X_13231_ _15063_/A VGND VGND VPWR VPWR _14529_/A sky130_fd_sc_hd__inv_2
X_10443_ _13522_/A _10442_/B _10442_/X _10360_/X VGND VGND VPWR VPWR _10443_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13162_ _13194_/A _13194_/B VGND VGND VPWR VPWR _13162_/Y sky130_fd_sc_hd__nor2_1
X_10374_ _10374_/A VGND VGND VPWR VPWR _11805_/A sky130_fd_sc_hd__inv_2
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12113_ _13906_/A _12149_/B VGND VGND VPWR VPWR _12210_/A sky130_fd_sc_hd__and2_1
XFILLER_123_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13093_ _13677_/A _13010_/B _13010_/Y VGND VGND VPWR VPWR _13093_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_104_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12044_ _13101_/A _11962_/B _11958_/A _11962_/B VGND VGND VPWR VPWR _12044_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15803_ _15673_/A _15673_/B _15673_/Y VGND VGND VPWR VPWR _15803_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15734_ _15752_/A _15734_/B VGND VGND VPWR VPWR _16112_/A sky130_fd_sc_hd__nor2_1
X_13995_ _13995_/A _13995_/B VGND VGND VPWR VPWR _13995_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12946_ _12946_/A VGND VGND VPWR VPWR _14944_/A sky130_fd_sc_hd__buf_1
X_15665_ _15665_/A _15665_/B VGND VGND VPWR VPWR _15665_/X sky130_fd_sc_hd__and2_1
XFILLER_73_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12877_ _12854_/A _12854_/B _12854_/Y VGND VGND VPWR VPWR _12877_/Y sky130_fd_sc_hd__o21ai_1
X_15596_ _16044_/A VGND VGND VPWR VPWR _15681_/A sky130_fd_sc_hd__inv_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14586_/A _14586_/B _14586_/Y VGND VGND VPWR VPWR _14616_/Y sky130_fd_sc_hd__o21ai_1
X_11828_ _11787_/A _11787_/B _11787_/Y VGND VGND VPWR VPWR _11828_/X sky130_fd_sc_hd__a21o_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14584_/A _14584_/B VGND VGND VPWR VPWR _14547_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11759_ _11759_/A _11759_/B VGND VGND VPWR VPWR _11759_/Y sky130_fd_sc_hd__nor2_1
X_14478_ _14477_/A _14477_/B _14477_/Y VGND VGND VPWR VPWR _14478_/X sky130_fd_sc_hd__a21o_1
X_16217_ _16217_/A VGND VGND VPWR VPWR _16217_/Y sky130_fd_sc_hd__inv_2
X_13429_ _13334_/A _13334_/B _13334_/A _13334_/B VGND VGND VPWR VPWR _13429_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16148_ _16148_/A VGND VGND VPWR VPWR _16148_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16079_ _16106_/A _16106_/B VGND VGND VPWR VPWR _16079_/X sky130_fd_sc_hd__and2_1
XFILLER_115_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08970_ _08970_/A _08970_/B VGND VGND VPWR VPWR _11389_/B sky130_fd_sc_hd__or2_1
XFILLER_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 wb_rst_i VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09522_ _09937_/A _09199_/Y _08703_/A _09199_/A VGND VGND VPWR VPWR _09522_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09453_ _09490_/A _09453_/B VGND VGND VPWR VPWR _09453_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08404_ _08361_/Y _08388_/Y _08404_/B1 _08388_/A _08419_/A VGND VGND VPWR VPWR _08653_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09384_ _09328_/A _09328_/B _09328_/X _09330_/A VGND VGND VPWR VPWR _11096_/A sky130_fd_sc_hd__a22o_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08335_ _08333_/Y _08334_/A _08333_/A _08334_/Y _08304_/A VGND VGND VPWR VPWR _09209_/B
+ sky130_fd_sc_hd__o221a_1
X_08266_ _08266_/A input13/X VGND VGND VPWR VPWR _08347_/A sky130_fd_sc_hd__nor2_1
XFILLER_106_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10090_ _10031_/X _10089_/X _10031_/X _10089_/X VGND VGND VPWR VPWR _10090_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12800_ _12778_/X _12799_/Y _12778_/X _12799_/Y VGND VGND VPWR VPWR _12854_/B sky130_fd_sc_hd__a2bb2o_1
X_13780_ _13778_/Y _13779_/Y _13716_/Y VGND VGND VPWR VPWR _13864_/A sky130_fd_sc_hd__o21ai_1
X_10992_ _12095_/A _11122_/B VGND VGND VPWR VPWR _10992_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _12717_/X _12730_/X _12717_/X _12730_/X VGND VGND VPWR VPWR _12781_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15450_ _15450_/A _15410_/X VGND VGND VPWR VPWR _15450_/X sky130_fd_sc_hd__or2b_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12662_/A VGND VGND VPWR VPWR _12662_/Y sky130_fd_sc_hd__inv_2
X_14401_ _15970_/A _14401_/B VGND VGND VPWR VPWR _14401_/X sky130_fd_sc_hd__or2_1
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11613_ _11612_/Y _11519_/X _11528_/X VGND VGND VPWR VPWR _11689_/A sky130_fd_sc_hd__o21ai_1
XFILLER_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12593_ _12619_/A _12619_/B VGND VGND VPWR VPWR _14226_/A sky130_fd_sc_hd__and2_1
X_15381_ _15381_/A _15337_/X VGND VGND VPWR VPWR _15381_/X sky130_fd_sc_hd__or2b_1
X_14332_ _14262_/A _14331_/Y _14262_/A _14331_/Y VGND VGND VPWR VPWR _14386_/A sky130_fd_sc_hd__a2bb2o_1
X_11544_ _13975_/A _11638_/B _11543_/Y VGND VGND VPWR VPWR _11544_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14263_ _15869_/A _14263_/B VGND VGND VPWR VPWR _14263_/Y sky130_fd_sc_hd__nand2_1
X_11475_ _11474_/A _11474_/B _11474_/Y _09393_/X VGND VGND VPWR VPWR _12440_/A sky130_fd_sc_hd__o211a_1
X_16002_ _16002_/A _15962_/X VGND VGND VPWR VPWR _16002_/X sky130_fd_sc_hd__or2b_1
X_13214_ _13205_/X _13213_/Y _13205_/X _13213_/Y VGND VGND VPWR VPWR _13306_/B sky130_fd_sc_hd__a2bb2o_1
X_10426_ _10426_/A _10426_/B VGND VGND VPWR VPWR _11792_/B sky130_fd_sc_hd__or2_1
X_14194_ _14113_/X _14193_/Y _14113_/X _14193_/Y VGND VGND VPWR VPWR _14195_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13145_ _15237_/A _13123_/B _13123_/Y VGND VGND VPWR VPWR _13145_/Y sky130_fd_sc_hd__o21ai_1
X_10357_ _12831_/A _10355_/B _10354_/X _10356_/Y VGND VGND VPWR VPWR _10357_/X sky130_fd_sc_hd__o22a_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _13019_/X _13075_/X _13019_/X _13075_/X VGND VGND VPWR VPWR _13111_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _12605_/A _10288_/B VGND VGND VPWR VPWR _10352_/A sky130_fd_sc_hd__or2_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12027_ _12055_/A VGND VGND VPWR VPWR _13190_/A sky130_fd_sc_hd__buf_1
XFILLER_66_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13978_ _13979_/A _13979_/B VGND VGND VPWR VPWR _13980_/A sky130_fd_sc_hd__and2_1
X_15717_ _15693_/Y _15716_/Y _15693_/Y _15716_/Y VGND VGND VPWR VPWR _15819_/B sky130_fd_sc_hd__a2bb2o_1
X_12929_ _12903_/Y _12927_/X _12928_/Y VGND VGND VPWR VPWR _12929_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15648_ _14377_/X _15647_/Y _14377_/X _15647_/Y VGND VGND VPWR VPWR _15667_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15579_ _15497_/X _15579_/B VGND VGND VPWR VPWR _15579_/X sky130_fd_sc_hd__and2b_1
XFILLER_115_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08953_ _08948_/Y _08951_/Y _08952_/Y VGND VGND VPWR VPWR _08960_/A sky130_fd_sc_hd__o21ai_1
XFILLER_130_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08884_ _08883_/Y _08865_/X _08883_/Y _08865_/X VGND VGND VPWR VPWR _08980_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09505_ _09505_/A VGND VGND VPWR VPWR _09505_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09436_/B VGND VGND VPWR VPWR _09436_/Y sky130_fd_sc_hd__nand2_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09367_ _09357_/X _09366_/X _09357_/X _09366_/X VGND VGND VPWR VPWR _09368_/A sky130_fd_sc_hd__a2bb2o_1
X_08318_ _08318_/A VGND VGND VPWR VPWR _08318_/Y sky130_fd_sc_hd__inv_2
X_09298_ _09298_/A _09298_/B VGND VGND VPWR VPWR _09299_/A sky130_fd_sc_hd__nand2_1
X_08249_ input3/X VGND VGND VPWR VPWR _08321_/A sky130_fd_sc_hd__inv_2
XFILLER_125_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11260_ _15446_/A _11188_/B _11188_/Y _11259_/X VGND VGND VPWR VPWR _11260_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10211_ _10463_/A _11711_/A VGND VGND VPWR VPWR _10281_/A sky130_fd_sc_hd__nand2_1
X_11191_ _09135_/Y _11190_/A _09135_/A _11190_/Y _09204_/X VGND VGND VPWR VPWR _13365_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_106_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10142_ _08770_/B _10132_/B _10133_/B VGND VGND VPWR VPWR _10143_/B sky130_fd_sc_hd__a21bo_1
X_14950_ _14935_/X _14949_/X _14935_/X _14949_/X VGND VGND VPWR VPWR _14976_/B sky130_fd_sc_hd__a2bb2o_1
X_10073_ _10073_/A _10073_/B VGND VGND VPWR VPWR _10073_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14881_ _14790_/A _14790_/B _14790_/A _14790_/B VGND VGND VPWR VPWR _14881_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13901_ _15414_/A _13956_/B VGND VGND VPWR VPWR _13901_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13832_ _14646_/A _13840_/B VGND VGND VPWR VPWR _13832_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13763_ _13763_/A _13763_/B VGND VGND VPWR VPWR _13763_/X sky130_fd_sc_hd__or2_1
X_15502_ _15481_/X _15501_/X _15481_/X _15501_/X VGND VGND VPWR VPWR _15544_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12714_ _12694_/A _12694_/B _12694_/Y _12713_/X VGND VGND VPWR VPWR _12714_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10975_ _10973_/A _10972_/Y _10973_/Y _10972_/A _11526_/A VGND VGND VPWR VPWR _11140_/B
+ sky130_fd_sc_hd__a221o_1
X_13694_ _13739_/A _13692_/X _13693_/X VGND VGND VPWR VPWR _13694_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12645_ _15554_/A VGND VGND VPWR VPWR _14984_/A sky130_fd_sc_hd__buf_1
X_15433_ _15433_/A _15563_/B VGND VGND VPWR VPWR _15433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12576_ _15524_/A VGND VGND VPWR VPWR _14910_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15364_ _15348_/X _15363_/X _15348_/X _15363_/X VGND VGND VPWR VPWR _15416_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14315_ _14335_/A _14315_/B VGND VGND VPWR VPWR _15962_/A sky130_fd_sc_hd__or2_1
X_11527_ _11612_/B VGND VGND VPWR VPWR _11528_/B sky130_fd_sc_hd__inv_2
XFILLER_129_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15295_ _15282_/X _15294_/Y _15282_/X _15294_/Y VGND VGND VPWR VPWR _15351_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14246_ _14362_/B VGND VGND VPWR VPWR _15778_/A sky130_fd_sc_hd__inv_2
X_11458_ _14132_/A _11363_/B _11363_/Y _12514_/A VGND VGND VPWR VPWR _12506_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14177_ _14278_/A VGND VGND VPWR VPWR _15906_/A sky130_fd_sc_hd__buf_1
X_10409_ _11780_/A _10409_/B VGND VGND VPWR VPWR _10409_/X sky130_fd_sc_hd__and2_1
X_11389_ _08912_/X _11389_/B VGND VGND VPWR VPWR _11389_/X sky130_fd_sc_hd__and2b_1
XFILLER_124_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13128_ _13037_/Y _13126_/X _13127_/Y VGND VGND VPWR VPWR _13128_/Y sky130_fd_sc_hd__o21ai_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13771_/A VGND VGND VPWR VPWR _15246_/A sky130_fd_sc_hd__buf_1
XFILLER_66_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09221_ _09221_/A _09221_/B VGND VGND VPWR VPWR _09802_/A sky130_fd_sc_hd__or2_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09152_ _09152_/A VGND VGND VPWR VPWR _09525_/B sky130_fd_sc_hd__inv_2
XFILLER_108_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09083_ _10013_/B _09076_/B _09077_/B VGND VGND VPWR VPWR _09766_/A sky130_fd_sc_hd__a21bo_1
XFILLER_1_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09985_ _09969_/Y _09983_/Y _09984_/Y VGND VGND VPWR VPWR _09987_/B sky130_fd_sc_hd__o21ai_1
X_08936_ _09503_/A _10103_/A _08935_/X VGND VGND VPWR VPWR _08936_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08867_ _09484_/A _08768_/Y _08770_/Y _08866_/X VGND VGND VPWR VPWR _08867_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08798_ _08798_/A VGND VGND VPWR VPWR _08798_/X sky130_fd_sc_hd__buf_1
XFILLER_72_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10760_ _11958_/A _10766_/B VGND VGND VPWR VPWR _10901_/A sky130_fd_sc_hd__and2_1
XFILLER_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10691_ _10809_/A _11990_/A VGND VGND VPWR VPWR _10691_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09419_ _10438_/A _09417_/Y _09418_/Y VGND VGND VPWR VPWR _09421_/B sky130_fd_sc_hd__o21ai_1
X_12430_ _12419_/A _12419_/B _12424_/X _12419_/Y _12429_/Y VGND VGND VPWR VPWR _12430_/X
+ sky130_fd_sc_hd__a32o_1
X_14100_ _14052_/X _14099_/X _14052_/X _14099_/X VGND VGND VPWR VPWR _14100_/Y sky130_fd_sc_hd__a2bb2oi_1
X_12361_ _12360_/Y _12253_/X _12287_/Y VGND VGND VPWR VPWR _12361_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12292_ _12250_/X _12291_/Y _12250_/X _12291_/Y VGND VGND VPWR VPWR _12294_/B sky130_fd_sc_hd__a2bb2o_1
X_15080_ _15029_/X _15079_/X _15029_/X _15079_/X VGND VGND VPWR VPWR _15081_/B sky130_fd_sc_hd__a2bb2o_1
X_11312_ _11312_/A _12179_/A VGND VGND VPWR VPWR _11312_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11243_ _11243_/A _11411_/B VGND VGND VPWR VPWR _14048_/A sky130_fd_sc_hd__or2_2
X_14031_ _13945_/X _14030_/Y _13945_/X _14030_/Y VGND VGND VPWR VPWR _14032_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11174_ _11103_/X _11173_/X _11103_/X _11173_/X VGND VGND VPWR VPWR _11176_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15982_ _15982_/A _15982_/B VGND VGND VPWR VPWR _15982_/X sky130_fd_sc_hd__or2_1
XFILLER_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10125_ _10125_/A _10125_/B VGND VGND VPWR VPWR _10126_/B sky130_fd_sc_hd__or2_1
XFILLER_121_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14933_ _14829_/X _14859_/A _14858_/X VGND VGND VPWR VPWR _14933_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10056_ _10055_/A _10055_/B _09954_/Y _10055_/X VGND VGND VPWR VPWR _10059_/A sky130_fd_sc_hd__a22o_1
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14864_ _14864_/A VGND VGND VPWR VPWR _15550_/A sky130_fd_sc_hd__buf_1
XFILLER_63_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14795_ _15458_/A VGND VGND VPWR VPWR _14798_/A sky130_fd_sc_hd__buf_1
X_13815_ _14619_/A _13850_/B VGND VGND VPWR VPWR _13815_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13746_ _13688_/X _13745_/Y _13688_/X _13745_/Y VGND VGND VPWR VPWR _13759_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10958_ _10081_/A _10956_/Y _09967_/Y _10956_/A _10957_/X VGND VGND VPWR VPWR _12078_/A
+ sky130_fd_sc_hd__o221a_1
X_16465_ _16357_/A _16465_/D VGND VGND VPWR VPWR _16465_/Q sky130_fd_sc_hd__dfxtp_1
X_13677_ _13677_/A VGND VGND VPWR VPWR _14501_/A sky130_fd_sc_hd__inv_2
XFILLER_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12628_ _14202_/A _12626_/X _12627_/X VGND VGND VPWR VPWR _12628_/X sky130_fd_sc_hd__o21a_1
X_15416_ _15416_/A _15416_/B VGND VGND VPWR VPWR _15416_/X sky130_fd_sc_hd__or2_1
X_10889_ _13088_/A _10747_/B _10747_/Y VGND VGND VPWR VPWR _10889_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16396_ _16396_/A _16396_/B _16396_/C _16457_/S VGND VGND VPWR VPWR _16397_/B sky130_fd_sc_hd__or4b_1
XFILLER_12_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12559_ _12559_/A VGND VGND VPWR VPWR _12559_/Y sky130_fd_sc_hd__inv_2
X_15347_ _15347_/A _15347_/B VGND VGND VPWR VPWR _15347_/X sky130_fd_sc_hd__or2_1
XFILLER_8_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15278_ _14584_/A _15252_/B _15252_/Y _15277_/X VGND VGND VPWR VPWR _15278_/X sky130_fd_sc_hd__a2bb2o_1
X_14229_ _14906_/A _14084_/B _14084_/X VGND VGND VPWR VPWR _14229_/X sky130_fd_sc_hd__o21ba_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09770_/A _09770_/B VGND VGND VPWR VPWR _09770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08721_ _08934_/A _08721_/B VGND VGND VPWR VPWR _09041_/A sky130_fd_sc_hd__nor2_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _08721_/B VGND VGND VPWR VPWR _08679_/A sky130_fd_sc_hd__buf_1
XFILLER_94_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08583_ _08714_/B VGND VGND VPWR VPWR _09467_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09204_ _11219_/B VGND VGND VPWR VPWR _09204_/X sky130_fd_sc_hd__buf_2
X_09135_ _09135_/A VGND VGND VPWR VPWR _09135_/Y sky130_fd_sc_hd__inv_2
X_09066_ _09066_/A VGND VGND VPWR VPWR _09829_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09968_ _10079_/A VGND VGND VPWR VPWR _09968_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08919_ _08919_/A VGND VGND VPWR VPWR _09541_/A sky130_fd_sc_hd__inv_2
XFILLER_94_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11930_ _11985_/B _11929_/Y _11985_/B _11929_/Y VGND VGND VPWR VPWR _11983_/B sky130_fd_sc_hd__o2bb2a_1
X_09899_ _09728_/A _09804_/Y _09857_/B VGND VGND VPWR VPWR _09899_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_85_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11861_ _11918_/B _11860_/X _11918_/B _11860_/X VGND VGND VPWR VPWR _11914_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14580_ _14580_/A _14580_/B VGND VGND VPWR VPWR _14580_/Y sky130_fd_sc_hd__nand2_1
X_11792_ _11792_/A _11792_/B VGND VGND VPWR VPWR _11792_/X sky130_fd_sc_hd__or2_1
XFILLER_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13600_ _13564_/A _13564_/B _13565_/A VGND VGND VPWR VPWR _13600_/Y sky130_fd_sc_hd__o21ai_1
X_10812_ _10811_/Y _10674_/X _10683_/Y VGND VGND VPWR VPWR _10812_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10743_ _11966_/A VGND VGND VPWR VPWR _13088_/A sky130_fd_sc_hd__buf_1
X_13531_ _12832_/A _12832_/B _10426_/B _12832_/Y VGND VGND VPWR VPWR _13531_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_53_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16250_ _16240_/Y _16248_/Y _16249_/Y VGND VGND VPWR VPWR _16250_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15201_ _15150_/X _15200_/Y _15150_/X _15200_/Y VGND VGND VPWR VPWR _15202_/B sky130_fd_sc_hd__a2bb2o_1
X_13462_ _11609_/Y _12677_/X _11691_/X VGND VGND VPWR VPWR _13462_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10674_ _10673_/Y _10555_/X _10564_/Y VGND VGND VPWR VPWR _10674_/X sky130_fd_sc_hd__o21a_1
X_16181_ _16189_/A _16181_/B VGND VGND VPWR VPWR _16262_/A sky130_fd_sc_hd__or2_1
X_13393_ _14114_/A _13438_/B VGND VGND VPWR VPWR _13393_/Y sky130_fd_sc_hd__nor2_1
X_12413_ _11611_/X _12422_/A _11611_/X _12422_/A VGND VGND VPWR VPWR _12426_/B sky130_fd_sc_hd__o2bb2a_1
X_12344_ _12344_/A _12344_/B VGND VGND VPWR VPWR _12344_/Y sky130_fd_sc_hd__nand2_1
X_15132_ _15075_/A _15075_/B _15075_/Y VGND VGND VPWR VPWR _15132_/Y sky130_fd_sc_hd__o21ai_1
X_15063_ _15063_/A _15063_/B VGND VGND VPWR VPWR _15063_/Y sky130_fd_sc_hd__nand2_1
X_14014_ _13955_/X _14013_/Y _13955_/X _14013_/Y VGND VGND VPWR VPWR _14060_/B sky130_fd_sc_hd__a2bb2o_1
X_12275_ _12373_/B _12274_/X _12373_/B _12274_/X VGND VGND VPWR VPWR _12370_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11226_ _13340_/A VGND VGND VPWR VPWR _12224_/A sky130_fd_sc_hd__inv_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11157_ _11312_/A _12266_/A VGND VGND VPWR VPWR _11157_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10108_ _10108_/A VGND VGND VPWR VPWR _10108_/Y sky130_fd_sc_hd__inv_2
X_15965_ _15999_/A _15963_/X _15964_/X VGND VGND VPWR VPWR _15966_/B sky130_fd_sc_hd__o21a_1
X_11088_ _11210_/A _11086_/X _11087_/X VGND VGND VPWR VPWR _11088_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15896_ _15896_/A _15896_/B VGND VGND VPWR VPWR _15896_/Y sky130_fd_sc_hd__nand2_1
X_14916_ _14916_/A _14916_/B VGND VGND VPWR VPWR _14916_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10039_ _10028_/X _10038_/Y _10028_/X _10038_/Y VGND VGND VPWR VPWR _10085_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14847_ _15178_/A _14848_/B VGND VGND VPWR VPWR _14849_/A sky130_fd_sc_hd__and2_1
XFILLER_17_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14778_ _14778_/A _14778_/B VGND VGND VPWR VPWR _14778_/X sky130_fd_sc_hd__and2_1
XFILLER_63_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13729_ _13771_/A _13771_/B VGND VGND VPWR VPWR _13807_/A sky130_fd_sc_hd__and2_1
X_16448_ _16446_/Y _16415_/X _16412_/Y _16429_/B _16447_/X VGND VGND VPWR VPWR _16448_/X
+ sky130_fd_sc_hd__o221a_1
X_16379_ _16317_/X _16378_/Y _16317_/X _16378_/Y VGND VGND VPWR VPWR _16396_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09822_ _09821_/A _09821_/B _09882_/B VGND VGND VPWR VPWR _09853_/A sky130_fd_sc_hd__a21bo_1
XFILLER_98_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09753_ _09997_/B VGND VGND VPWR VPWR _09753_/Y sky130_fd_sc_hd__inv_2
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ _09937_/A _08704_/B VGND VGND VPWR VPWR _09342_/A sky130_fd_sc_hd__or2_1
XFILLER_67_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09684_ _09684_/A _09684_/B VGND VGND VPWR VPWR _09687_/B sky130_fd_sc_hd__or2_1
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08635_ _08635_/A VGND VGND VPWR VPWR _10111_/B sky130_fd_sc_hd__inv_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08566_ _09858_/A VGND VGND VPWR VPWR _09734_/A sky130_fd_sc_hd__inv_2
XFILLER_23_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08497_ _08298_/X _08496_/X _08298_/X _08496_/X VGND VGND VPWR VPWR _08660_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09118_ _09705_/A _09118_/B VGND VGND VPWR VPWR _09118_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10390_ _13522_/A _10442_/B _13522_/A _10442_/B VGND VGND VPWR VPWR _10390_/X sky130_fd_sc_hd__a2bb2o_1
X_09049_ _08713_/A _08713_/B _08713_/X _09048_/Y VGND VGND VPWR VPWR _09050_/A sky130_fd_sc_hd__a22o_1
XFILLER_2_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12060_ _12022_/Y _12058_/X _12059_/Y VGND VGND VPWR VPWR _12060_/X sky130_fd_sc_hd__o21a_1
X_11011_ _11011_/A _10922_/X VGND VGND VPWR VPWR _11011_/X sky130_fd_sc_hd__or2b_1
XFILLER_2_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15750_ _14914_/A _14914_/B _14914_/Y VGND VGND VPWR VPWR _15750_/X sky130_fd_sc_hd__o21a_1
X_12962_ _13720_/A VGND VGND VPWR VPWR _14669_/A sky130_fd_sc_hd__inv_2
XFILLER_58_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15681_ _15681_/A _15681_/B VGND VGND VPWR VPWR _15681_/Y sky130_fd_sc_hd__nand2_1
X_14701_ _14655_/X _14700_/Y _14655_/X _14700_/Y VGND VGND VPWR VPWR _14733_/B sky130_fd_sc_hd__a2bb2o_1
X_12893_ _12846_/A _12846_/B _12846_/Y VGND VGND VPWR VPWR _12893_/Y sky130_fd_sc_hd__o21ai_1
X_11913_ _11913_/A _11913_/B VGND VGND VPWR VPWR _11913_/X sky130_fd_sc_hd__or2_1
XFILLER_18_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14632_ _14578_/A _14578_/B _14578_/Y VGND VGND VPWR VPWR _14632_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11844_ _11818_/Y _11842_/X _11843_/Y VGND VGND VPWR VPWR _11844_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14576_/A _14576_/B VGND VGND VPWR VPWR _14563_/Y sky130_fd_sc_hd__nor2_1
X_11775_ _11775_/A _11775_/B VGND VGND VPWR VPWR _11775_/X sky130_fd_sc_hd__and2_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16324_/A _16324_/B VGND VGND VPWR VPWR _16302_/Y sky130_fd_sc_hd__nor2_1
X_14494_ _14463_/A _14463_/B _14463_/Y VGND VGND VPWR VPWR _14494_/Y sky130_fd_sc_hd__o21ai_1
X_10726_ _11901_/A VGND VGND VPWR VPWR _13693_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13514_ _13516_/A VGND VGND VPWR VPWR _15038_/A sky130_fd_sc_hd__buf_1
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16233_ _16233_/A VGND VGND VPWR VPWR _16233_/Y sky130_fd_sc_hd__inv_2
X_13445_ _13384_/Y _13443_/X _13444_/Y VGND VGND VPWR VPWR _13445_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10657_ _11021_/A _10657_/B VGND VGND VPWR VPWR _10657_/X sky130_fd_sc_hd__and2_1
XFILLER_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16164_ _16111_/X _16163_/X _16111_/X _16163_/X VGND VGND VPWR VPWR _16165_/B sky130_fd_sc_hd__a2bb2oi_1
X_13376_ _13313_/A _13313_/B _13313_/A _13313_/B VGND VGND VPWR VPWR _13376_/X sky130_fd_sc_hd__a2bb2o_1
X_10588_ _11904_/A _10641_/B VGND VGND VPWR VPWR _10588_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16095_ _16091_/Y _16213_/A _16094_/Y VGND VGND VPWR VPWR _16099_/B sky130_fd_sc_hd__o21ai_1
XFILLER_126_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12327_ _12227_/A _12227_/B _12227_/Y VGND VGND VPWR VPWR _12327_/Y sky130_fd_sc_hd__o21ai_1
X_15115_ _15097_/X _15114_/Y _15097_/X _15114_/Y VGND VGND VPWR VPWR _15116_/B sky130_fd_sc_hd__a2bb2o_1
X_12258_ _12257_/Y _12164_/X _12187_/Y VGND VGND VPWR VPWR _12258_/X sky130_fd_sc_hd__o21a_1
X_15046_ _15046_/A _15046_/B VGND VGND VPWR VPWR _15046_/X sky130_fd_sc_hd__or2_1
X_11209_ _12215_/A VGND VGND VPWR VPWR _11449_/A sky130_fd_sc_hd__buf_1
XFILLER_79_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12189_ _12164_/X _12188_/Y _12164_/X _12188_/Y VGND VGND VPWR VPWR _12254_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15948_ _15948_/A _15948_/B VGND VGND VPWR VPWR _15948_/X sky130_fd_sc_hd__or2_1
XFILLER_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15879_ _14226_/X _15841_/X _14226_/X _15841_/X VGND VGND VPWR VPWR _15888_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08420_ _08418_/A _08343_/Y _08418_/Y _08343_/A _08441_/A VGND VGND VPWR VPWR _09217_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08351_ _09221_/B VGND VGND VPWR VPWR _08351_/Y sky130_fd_sc_hd__inv_2
X_08282_ _08282_/A VGND VGND VPWR VPWR _08399_/B sky130_fd_sc_hd__inv_2
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09805_ _09803_/A _09803_/B _09804_/Y VGND VGND VPWR VPWR _09855_/B sky130_fd_sc_hd__a21oi_1
X_09736_ _09736_/A _09736_/B VGND VGND VPWR VPWR _09739_/A sky130_fd_sc_hd__or2_1
XFILLER_55_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09667_ _09574_/Y _09665_/X _09666_/Y VGND VGND VPWR VPWR _09667_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_131_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08618_ _09456_/A _09221_/B _10016_/A _08351_/Y VGND VGND VPWR VPWR _08618_/X sky130_fd_sc_hd__o22a_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09598_ _08795_/X _09492_/B _09492_/Y VGND VGND VPWR VPWR _09598_/X sky130_fd_sc_hd__a21o_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08549_/A VGND VGND VPWR VPWR _08549_/Y sky130_fd_sc_hd__inv_2
X_11560_ _11472_/X _11559_/X _11472_/X _11559_/X VGND VGND VPWR VPWR _11561_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10511_ _11835_/A VGND VGND VPWR VPWR _15143_/A sky130_fd_sc_hd__buf_1
XFILLER_50_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13230_ _14739_/A _13297_/B VGND VGND VPWR VPWR _13230_/Y sky130_fd_sc_hd__nor2_1
X_11491_ _12362_/A _11491_/B VGND VGND VPWR VPWR _11491_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10442_ _11755_/A _10442_/B VGND VGND VPWR VPWR _10442_/X sky130_fd_sc_hd__and2_1
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13161_ _13112_/X _13160_/Y _13112_/X _13160_/Y VGND VGND VPWR VPWR _13194_/B sky130_fd_sc_hd__a2bb2o_1
X_10373_ _10455_/A _11219_/A VGND VGND VPWR VPWR _10374_/A sky130_fd_sc_hd__or2_1
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13092_ _15264_/A _13105_/B VGND VGND VPWR VPWR _13092_/Y sky130_fd_sc_hd__nor2_1
X_12112_ _12060_/X _12111_/Y _12060_/X _12111_/Y VGND VGND VPWR VPWR _12149_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_97_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12043_ _12043_/A VGND VGND VPWR VPWR _12043_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15802_ _16104_/A _15805_/B VGND VGND VPWR VPWR _15802_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15733_ _14919_/X _15732_/X _14919_/X _15732_/X VGND VGND VPWR VPWR _15734_/B sky130_fd_sc_hd__a2bb2oi_1
X_13994_ _15422_/A _13995_/B VGND VGND VPWR VPWR _13994_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12945_ _12871_/Y _12943_/X _12944_/Y VGND VGND VPWR VPWR _12945_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15664_ _15665_/A _15665_/B VGND VGND VPWR VPWR _15775_/B sky130_fd_sc_hd__or2_1
X_12876_ _12940_/A VGND VGND VPWR VPWR _14600_/A sky130_fd_sc_hd__buf_1
X_15595_ _15595_/A _15595_/B VGND VGND VPWR VPWR _16044_/A sky130_fd_sc_hd__or2_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _14615_/A VGND VGND VPWR VPWR _15343_/A sky130_fd_sc_hd__buf_1
X_11827_ _13606_/A _11837_/B VGND VGND VPWR VPWR _11827_/Y sky130_fd_sc_hd__nor2_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _14519_/X _14545_/X _14519_/X _14545_/X VGND VGND VPWR VPWR _14584_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11758_ _11757_/A _11757_/B _11757_/X _11750_/B VGND VGND VPWR VPWR _11803_/B sky130_fd_sc_hd__a22o_1
XFILLER_119_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10709_ _11907_/A VGND VGND VPWR VPWR _13697_/A sky130_fd_sc_hd__buf_1
X_14477_ _14477_/A _14477_/B VGND VGND VPWR VPWR _14477_/Y sky130_fd_sc_hd__nor2_1
X_11689_ _11689_/A VGND VGND VPWR VPWR _11689_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16216_ _16099_/A _15800_/B _15800_/Y VGND VGND VPWR VPWR _16218_/A sky130_fd_sc_hd__o21ai_1
X_13428_ _14106_/A _13431_/B VGND VGND VPWR VPWR _13428_/Y sky130_fd_sc_hd__nor2_1
X_16147_ _16147_/A VGND VGND VPWR VPWR _16147_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13359_ _13340_/A _13340_/B _13340_/X _13358_/X VGND VGND VPWR VPWR _13359_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16078_ _16037_/X _16077_/Y _16037_/X _16077_/Y VGND VGND VPWR VPWR _16106_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15029_ _15082_/A _15027_/X _15028_/X VGND VGND VPWR VPWR _15029_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 wbs_adr_i[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09521_ _09519_/Y _09520_/X _09519_/Y _09520_/X VGND VGND VPWR VPWR _09521_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_64_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09452_ _09452_/A _09531_/A VGND VGND VPWR VPWR _09452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08403_ _08852_/A _08398_/Y _08402_/X VGND VGND VPWR VPWR _08403_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09383_ _09432_/B _09383_/B VGND VGND VPWR VPWR _09383_/X sky130_fd_sc_hd__or2_1
X_08334_ _08334_/A VGND VGND VPWR VPWR _08334_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08265_ input29/X VGND VGND VPWR VPWR _08266_/A sky130_fd_sc_hd__inv_2
XFILLER_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10991_ _10952_/X _10990_/X _10952_/X _10990_/X VGND VGND VPWR VPWR _11122_/B sky130_fd_sc_hd__a2bb2o_1
X_09719_ _09720_/A _09720_/B VGND VGND VPWR VPWR _09719_/Y sky130_fd_sc_hd__nor2_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12730_ _12686_/A _12686_/B _12686_/Y VGND VGND VPWR VPWR _12730_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _10453_/Y _12660_/Y _10379_/Y VGND VGND VPWR VPWR _12662_/A sky130_fd_sc_hd__o21ai_1
X_14400_ _14285_/X _14399_/X _14285_/X _14399_/X VGND VGND VPWR VPWR _14400_/Y sky130_fd_sc_hd__a2bb2oi_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11612_ _11612_/A _11612_/B VGND VGND VPWR VPWR _11612_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12592_ _12589_/Y _12591_/Y _12589_/A _12591_/A _12500_/A VGND VGND VPWR VPWR _12619_/B
+ sky130_fd_sc_hd__o221a_1
X_15380_ _15406_/A _15406_/B VGND VGND VPWR VPWR _15456_/A sky130_fd_sc_hd__and2_1
XFILLER_11_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14331_ _15869_/A _14263_/B _14263_/Y VGND VGND VPWR VPWR _14331_/Y sky130_fd_sc_hd__o21ai_1
X_11543_ _12387_/A _11638_/B VGND VGND VPWR VPWR _11543_/Y sky130_fd_sc_hd__nand2_1
X_14262_ _14262_/A VGND VGND VPWR VPWR _14262_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11474_ _11474_/A _11474_/B VGND VGND VPWR VPWR _11474_/Y sky130_fd_sc_hd__nand2_1
X_16001_ _16046_/A _16046_/B VGND VGND VPWR VPWR _16001_/Y sky130_fd_sc_hd__nor2_1
X_14193_ _13438_/A _14115_/A _14079_/Y VGND VGND VPWR VPWR _14193_/Y sky130_fd_sc_hd__a21oi_1
X_13213_ _13206_/A _13206_/B _13206_/Y VGND VGND VPWR VPWR _13213_/Y sky130_fd_sc_hd__o21ai_1
X_10425_ _10425_/A VGND VGND VPWR VPWR _10426_/B sky130_fd_sc_hd__inv_2
XFILLER_124_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13144_ _13206_/A _13206_/B VGND VGND VPWR VPWR _13144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10356_ _10356_/A VGND VGND VPWR VPWR _10356_/Y sky130_fd_sc_hd__inv_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13075_ _13075_/A _13020_/X VGND VGND VPWR VPWR _13075_/X sky130_fd_sc_hd__or2b_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _10287_/A VGND VGND VPWR VPWR _12605_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12026_ _13192_/A _12057_/B VGND VGND VPWR VPWR _12026_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13977_ _13974_/X _13998_/A _13974_/X _13998_/A VGND VGND VPWR VPWR _13979_/B sky130_fd_sc_hd__a2bb2o_1
X_15716_ _15694_/A _15694_/B _15694_/Y VGND VGND VPWR VPWR _15716_/Y sky130_fd_sc_hd__o21ai_1
X_12928_ _12928_/A _12928_/B VGND VGND VPWR VPWR _12928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15647_ _14378_/A _14378_/B _14378_/Y VGND VGND VPWR VPWR _15647_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12859_ _12795_/Y _12857_/X _12858_/Y VGND VGND VPWR VPWR _12859_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15578_ _16055_/A _15696_/B VGND VGND VPWR VPWR _15578_/Y sky130_fd_sc_hd__nor2_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14529_ _14529_/A _14529_/B VGND VGND VPWR VPWR _14529_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08952_ _08952_/A _08952_/B VGND VGND VPWR VPWR _08952_/Y sky130_fd_sc_hd__nand2_1
X_08883_ _08778_/A _08778_/B _08778_/Y VGND VGND VPWR VPWR _08883_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09504_ _08847_/A _09460_/A _09826_/B _09460_/Y VGND VGND VPWR VPWR _09505_/A sky130_fd_sc_hd__o22a_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09435_ _09763_/A _09436_/B VGND VGND VPWR VPWR _09435_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09366_ _09476_/B _09862_/A _09349_/A VGND VGND VPWR VPWR _09366_/X sky130_fd_sc_hd__o21a_1
X_09297_ _09297_/A VGND VGND VPWR VPWR _09297_/Y sky130_fd_sc_hd__inv_2
X_08317_ _08317_/A _08317_/B VGND VGND VPWR VPWR _08318_/A sky130_fd_sc_hd__or2_1
X_08248_ input4/X _08248_/B VGND VGND VPWR VPWR _08317_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10210_ _10210_/A VGND VGND VPWR VPWR _11711_/A sky130_fd_sc_hd__inv_2
XFILLER_106_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11190_ _11190_/A VGND VGND VPWR VPWR _11190_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10141_ _10143_/A VGND VGND VPWR VPWR _10239_/B sky130_fd_sc_hd__buf_1
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10072_ _10071_/A _10071_/B _09970_/A _10071_/X VGND VGND VPWR VPWR _10075_/A sky130_fd_sc_hd__a22o_1
X_13900_ _13855_/X _13899_/Y _13855_/X _13899_/Y VGND VGND VPWR VPWR _13956_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14880_ _14880_/A VGND VGND VPWR VPWR _15542_/A sky130_fd_sc_hd__buf_1
X_13831_ _13756_/X _13830_/Y _13756_/X _13830_/Y VGND VGND VPWR VPWR _13840_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13762_ _13822_/A _13760_/X _13761_/X VGND VGND VPWR VPWR _13762_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10974_ _10974_/A VGND VGND VPWR VPWR _11526_/A sky130_fd_sc_hd__clkbuf_2
X_15501_ _15449_/A _15449_/B _15449_/A _15449_/B VGND VGND VPWR VPWR _15501_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12713_ _12696_/A _12696_/B _12696_/Y _12712_/X VGND VGND VPWR VPWR _12713_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13693_ _13693_/A _13693_/B VGND VGND VPWR VPWR _13693_/X sky130_fd_sc_hd__or2_1
XFILLER_43_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12644_ _12643_/A _12643_/B _12643_/Y _11707_/X VGND VGND VPWR VPWR _12650_/A sky130_fd_sc_hd__o211ai_1
X_15432_ _15421_/Y _15431_/Y _15421_/Y _15431_/Y VGND VGND VPWR VPWR _15563_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12575_ _12575_/A VGND VGND VPWR VPWR _15524_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15363_ _15363_/A _15349_/X VGND VGND VPWR VPWR _15363_/X sky130_fd_sc_hd__or2b_1
XFILLER_11_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14314_ _13439_/X _14313_/X _13439_/X _14313_/X VGND VGND VPWR VPWR _14315_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11526_ _11526_/A _11526_/B VGND VGND VPWR VPWR _11612_/B sky130_fd_sc_hd__or2_1
X_15294_ _15237_/A _15237_/B _15237_/Y VGND VGND VPWR VPWR _15294_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14245_ _14245_/A _14362_/B VGND VGND VPWR VPWR _14248_/A sky130_fd_sc_hd__or2_1
X_11457_ _14126_/A _11370_/B _11370_/Y _12522_/A VGND VGND VPWR VPWR _12514_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14176_ _14282_/A _14176_/B VGND VGND VPWR VPWR _14278_/A sky130_fd_sc_hd__or2_1
X_11388_ _14108_/A VGND VGND VPWR VPWR _12349_/A sky130_fd_sc_hd__inv_2
X_10408_ _10358_/X _10407_/X _10358_/X _10407_/X VGND VGND VPWR VPWR _10409_/B sky130_fd_sc_hd__a2bb2o_1
X_13127_ _13985_/A _13127_/B VGND VGND VPWR VPWR _13127_/Y sky130_fd_sc_hd__nand2_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _09707_/A _09707_/B _09707_/Y VGND VGND VPWR VPWR _10339_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_100_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13058_ _13058_/A VGND VGND VPWR VPWR _13771_/A sky130_fd_sc_hd__inv_2
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12009_ _13701_/A _12068_/B _12008_/Y VGND VGND VPWR VPWR _12009_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09220_ _09220_/A VGND VGND VPWR VPWR _09220_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09151_ _09518_/A _09148_/X _09148_/X _08524_/Y VGND VGND VPWR VPWR _09152_/A sky130_fd_sc_hd__o2bb2a_1
X_09082_ _09763_/A VGND VGND VPWR VPWR _09436_/A sky130_fd_sc_hd__buf_1
XFILLER_30_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09984_ _09984_/A _09984_/B VGND VGND VPWR VPWR _09984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08935_ _08935_/A _08935_/B VGND VGND VPWR VPWR _08935_/X sky130_fd_sc_hd__or2_1
XFILLER_57_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08866_ _09486_/A _08776_/Y _08778_/Y _08865_/X VGND VGND VPWR VPWR _08866_/X sky130_fd_sc_hd__o22a_1
XFILLER_72_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08797_ _08797_/A VGND VGND VPWR VPWR _08798_/A sky130_fd_sc_hd__inv_2
XFILLER_84_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10690_ _11990_/A VGND VGND VPWR VPWR _12692_/A sky130_fd_sc_hd__buf_1
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09418_ _09418_/A _09418_/B VGND VGND VPWR VPWR _09418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09349_ _09349_/A VGND VGND VPWR VPWR _09349_/Y sky130_fd_sc_hd__inv_2
X_12360_ _12360_/A _12360_/B VGND VGND VPWR VPWR _12360_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11311_ _12266_/A VGND VGND VPWR VPWR _12179_/A sky130_fd_sc_hd__inv_2
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12291_ _13204_/A _12358_/B _12290_/Y VGND VGND VPWR VPWR _12291_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11242_ _12230_/A _11242_/B VGND VGND VPWR VPWR _11242_/Y sky130_fd_sc_hd__nand2_1
X_14030_ _15404_/A _13946_/B _13946_/Y VGND VGND VPWR VPWR _14030_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11173_ _14664_/A _11276_/B _11276_/A _11276_/B VGND VGND VPWR VPWR _11173_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10124_ _10124_/A _10124_/B VGND VGND VPWR VPWR _10125_/B sky130_fd_sc_hd__or2_1
X_15981_ _15982_/A _15982_/B VGND VGND VPWR VPWR _15988_/A sky130_fd_sc_hd__and2_1
XFILLER_94_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14932_ _15433_/A VGND VGND VPWR VPWR _15563_/A sky130_fd_sc_hd__buf_1
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10055_ _10055_/A _10055_/B VGND VGND VPWR VPWR _10055_/X sky130_fd_sc_hd__or2_1
X_14863_ _15552_/A _14928_/B VGND VGND VPWR VPWR _14863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13814_ _13766_/X _13813_/X _13766_/X _13813_/X VGND VGND VPWR VPWR _13850_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14794_ _14794_/A _14794_/B VGND VGND VPWR VPWR _14794_/X sky130_fd_sc_hd__and2_1
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13745_ _14497_/A _13689_/B _13689_/Y VGND VGND VPWR VPWR _13745_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10957_ _10957_/A VGND VGND VPWR VPWR _10957_/X sky130_fd_sc_hd__clkbuf_2
X_16464_ _16357_/A _16464_/D VGND VGND VPWR VPWR _16464_/Q sky130_fd_sc_hd__dfxtp_1
X_13676_ _14497_/A _13689_/B VGND VGND VPWR VPWR _13676_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12627_ _12627_/A _12627_/B VGND VGND VPWR VPWR _12627_/X sky130_fd_sc_hd__or2_1
X_15415_ _15444_/A _15413_/X _15414_/X VGND VGND VPWR VPWR _15415_/X sky130_fd_sc_hd__o21a_1
X_10888_ _12037_/A VGND VGND VPWR VPWR _13825_/A sky130_fd_sc_hd__buf_1
X_16395_ _16395_/A VGND VGND VPWR VPWR _16396_/B sky130_fd_sc_hd__inv_2
X_12558_ _12554_/Y _12557_/Y _12554_/A _12557_/A _11707_/A VGND VGND VPWR VPWR _12625_/A
+ sky130_fd_sc_hd__o221a_1
X_15346_ _15369_/A _15344_/X _15345_/X VGND VGND VPWR VPWR _15346_/X sky130_fd_sc_hd__o21a_1
X_12489_ _12479_/Y _12488_/X _12479_/Y _12488_/X VGND VGND VPWR VPWR _12489_/X sky130_fd_sc_hd__a2bb2o_1
X_15277_ _14582_/A _15255_/B _15255_/Y _15276_/X VGND VGND VPWR VPWR _15277_/X sky130_fd_sc_hd__a2bb2o_1
X_11509_ _09964_/X _11509_/B VGND VGND VPWR VPWR _11510_/B sky130_fd_sc_hd__and2b_1
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14228_ _15878_/A _14254_/B VGND VGND VPWR VPWR _14228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14159_ _14207_/A VGND VGND VPWR VPWR _14282_/A sky130_fd_sc_hd__buf_1
XFILLER_112_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _08856_/B VGND VGND VPWR VPWR _09540_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08651_ _08856_/B VGND VGND VPWR VPWR _08721_/B sky130_fd_sc_hd__inv_2
XFILLER_94_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08582_ _09454_/B VGND VGND VPWR VPWR _08714_/B sky130_fd_sc_hd__inv_2
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09203_ _11249_/B VGND VGND VPWR VPWR _11219_/B sky130_fd_sc_hd__buf_2
X_09134_ _09555_/B _09036_/B _09037_/B VGND VGND VPWR VPWR _09135_/A sky130_fd_sc_hd__a21bo_1
XFILLER_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09065_ _09503_/B _09064_/A _09826_/B _09064_/Y VGND VGND VPWR VPWR _09069_/A sky130_fd_sc_hd__o22a_1
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09967_ _10081_/A VGND VGND VPWR VPWR _09967_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08918_ _09677_/A VGND VGND VPWR VPWR _08930_/A sky130_fd_sc_hd__inv_2
XFILLER_57_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09898_/A _09898_/B VGND VGND VPWR VPWR _09901_/A sky130_fd_sc_hd__and2_1
XFILLER_18_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08849_ _08935_/B VGND VGND VPWR VPWR _10103_/A sky130_fd_sc_hd__inv_2
XFILLER_72_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11860_ _11860_/A _11859_/X VGND VGND VPWR VPWR _11860_/X sky130_fd_sc_hd__or2b_1
X_11791_ _11791_/A _11791_/B VGND VGND VPWR VPWR _11791_/X sky130_fd_sc_hd__and2_1
XFILLER_41_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10811_ _11992_/A _10811_/B VGND VGND VPWR VPWR _10811_/Y sky130_fd_sc_hd__nor2_1
X_13530_ _13530_/A _13530_/B VGND VGND VPWR VPWR _13530_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10742_ _10740_/A _10741_/A _10740_/Y _10741_/Y _09672_/A VGND VGND VPWR VPWR _11966_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_41_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15200_ _15134_/A _15134_/B _15134_/Y VGND VGND VPWR VPWR _15200_/Y sky130_fd_sc_hd__o21ai_1
X_13461_ _15425_/A _12863_/B _12863_/Y _12948_/X VGND VGND VPWR VPWR _13461_/Y sky130_fd_sc_hd__o2bb2ai_1
X_10673_ _11920_/A _10673_/B VGND VGND VPWR VPWR _10673_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16180_ _16107_/X _16179_/X _16107_/X _16179_/X VGND VGND VPWR VPWR _16181_/B sky130_fd_sc_hd__a2bb2oi_1
X_13392_ _13362_/X _13391_/X _13362_/X _13391_/X VGND VGND VPWR VPWR _13438_/B sky130_fd_sc_hd__a2bb2o_1
X_12412_ _11612_/A _11528_/B _12376_/X VGND VGND VPWR VPWR _12422_/A sky130_fd_sc_hd__o21ai_1
X_12343_ _12241_/X _12342_/Y _12241_/X _12342_/Y VGND VGND VPWR VPWR _12559_/A sky130_fd_sc_hd__a2bb2o_1
X_15131_ _15131_/A _15131_/B VGND VGND VPWR VPWR _15131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15062_ _15041_/X _15061_/X _15041_/X _15061_/X VGND VGND VPWR VPWR _15063_/B sky130_fd_sc_hd__a2bb2o_1
X_12274_ _12274_/A _12273_/X VGND VGND VPWR VPWR _12274_/X sky130_fd_sc_hd__or2b_1
XFILLER_5_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11225_ _11225_/A _11249_/B VGND VGND VPWR VPWR _13340_/A sky130_fd_sc_hd__or2_1
X_14013_ _15414_/A _13956_/B _13956_/Y VGND VGND VPWR VPWR _14013_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11156_ _11155_/A _11155_/B _11155_/Y _10982_/X VGND VGND VPWR VPWR _12266_/A sky130_fd_sc_hd__o211a_1
XFILLER_122_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15964_ _15964_/A _15964_/B VGND VGND VPWR VPWR _15964_/X sky130_fd_sc_hd__or2_1
X_11087_ _13910_/A _11087_/B VGND VGND VPWR VPWR _11087_/X sky130_fd_sc_hd__or2_1
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10107_ _10177_/A _10177_/B _10106_/Y VGND VGND VPWR VPWR _10109_/A sky130_fd_sc_hd__o21ai_1
X_14915_ _14889_/Y _14913_/X _14914_/Y VGND VGND VPWR VPWR _14915_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10038_ _10038_/A _10038_/B VGND VGND VPWR VPWR _10038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15895_ _15871_/Y _15893_/X _15894_/Y VGND VGND VPWR VPWR _15895_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14846_ _14837_/X _14845_/Y _14837_/X _14845_/Y VGND VGND VPWR VPWR _14848_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14777_ _14740_/X _14776_/X _14740_/X _14776_/X VGND VGND VPWR VPWR _14778_/B sky130_fd_sc_hd__a2bb2o_1
X_13728_ _13700_/X _13727_/X _13700_/X _13727_/X VGND VGND VPWR VPWR _13771_/B sky130_fd_sc_hd__a2bb2o_1
X_11989_ _12075_/A VGND VGND VPWR VPWR _12777_/A sky130_fd_sc_hd__buf_1
XFILLER_44_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16447_ _16447_/A _16447_/B VGND VGND VPWR VPWR _16447_/X sky130_fd_sc_hd__or2_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13659_ _15125_/A _13638_/B _13638_/Y VGND VGND VPWR VPWR _13659_/Y sky130_fd_sc_hd__o21ai_1
X_16378_ _16378_/A1 _16318_/B _16318_/Y VGND VGND VPWR VPWR _16378_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15329_ _15329_/A _15329_/B VGND VGND VPWR VPWR _15329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09821_ _09821_/A _09821_/B VGND VGND VPWR VPWR _09882_/B sky130_fd_sc_hd__or2_1
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09752_ _10087_/A VGND VGND VPWR VPWR _09997_/B sky130_fd_sc_hd__buf_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _08703_/A VGND VGND VPWR VPWR _09937_/A sky130_fd_sc_hd__inv_2
XFILLER_104_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09683_ _09683_/A _09683_/B VGND VGND VPWR VPWR _09686_/A sky130_fd_sc_hd__or2_1
XFILLER_27_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08634_ _08634_/A VGND VGND VPWR VPWR _09462_/B sky130_fd_sc_hd__inv_2
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08565_ _10012_/A _08565_/B VGND VGND VPWR VPWR _09858_/A sky130_fd_sc_hd__or2_2
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08496_ _08239_/Y _08699_/A _08237_/A _08235_/B VGND VGND VPWR VPWR _08496_/X sky130_fd_sc_hd__o22a_2
XFILLER_23_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09117_ _09117_/A VGND VGND VPWR VPWR _09117_/Y sky130_fd_sc_hd__inv_2
X_09048_ _08714_/Y _09047_/Y _08730_/X VGND VGND VPWR VPWR _09048_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11010_ _15063_/A VGND VGND VPWR VPWR _13902_/A sky130_fd_sc_hd__buf_1
XFILLER_104_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12961_ _14749_/A _13032_/B VGND VGND VPWR VPWR _13045_/A sky130_fd_sc_hd__and2_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15680_ _15607_/Y _15678_/X _15679_/Y VGND VGND VPWR VPWR _15680_/X sky130_fd_sc_hd__o21a_1
X_14700_ _15341_/A _14656_/B _14656_/Y VGND VGND VPWR VPWR _14700_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12892_ _12932_/A VGND VGND VPWR VPWR _14467_/A sky130_fd_sc_hd__buf_1
X_11912_ _13552_/A _11911_/B _11911_/X _11846_/X VGND VGND VPWR VPWR _11912_/X sky130_fd_sc_hd__o22a_1
XFILLER_18_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14631_ _14631_/A VGND VGND VPWR VPWR _15335_/A sky130_fd_sc_hd__buf_1
X_11843_ _11843_/A _11843_/B VGND VGND VPWR VPWR _11843_/Y sky130_fd_sc_hd__nand2_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16256_/X _16300_/Y _16256_/X _16300_/Y VGND VGND VPWR VPWR _16324_/B sky130_fd_sc_hd__o2bb2a_1
X_14562_ _14511_/X _14561_/X _14511_/X _14561_/X VGND VGND VPWR VPWR _14576_/B sky130_fd_sc_hd__a2bb2o_1
X_11774_ _11741_/B _11773_/Y _11741_/B _11773_/Y VGND VGND VPWR VPWR _11775_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _14493_/A VGND VGND VPWR VPWR _15205_/A sky130_fd_sc_hd__buf_1
X_10725_ _11970_/A VGND VGND VPWR VPWR _13078_/A sky130_fd_sc_hd__buf_1
X_13513_ _13513_/A _13513_/B VGND VGND VPWR VPWR _13513_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16232_ _16084_/A _16084_/B _16084_/Y VGND VGND VPWR VPWR _16234_/A sky130_fd_sc_hd__o21ai_1
X_13444_ _13444_/A _13444_/B VGND VGND VPWR VPWR _13444_/Y sky130_fd_sc_hd__nand2_1
X_10656_ _12936_/A VGND VGND VPWR VPWR _11933_/A sky130_fd_sc_hd__inv_2
XFILLER_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16163_ _16070_/X _16163_/B VGND VGND VPWR VPWR _16163_/X sky130_fd_sc_hd__and2b_1
X_13375_ _13450_/A _13450_/B VGND VGND VPWR VPWR _13375_/Y sky130_fd_sc_hd__nor2_1
X_10587_ _10532_/X _10586_/Y _10532_/X _10586_/Y VGND VGND VPWR VPWR _10641_/B sky130_fd_sc_hd__a2bb2o_1
X_15114_ _15057_/A _15057_/B _15057_/Y VGND VGND VPWR VPWR _15114_/Y sky130_fd_sc_hd__o21ai_1
X_16094_ _16094_/A _16094_/B VGND VGND VPWR VPWR _16094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12326_ _12329_/A _12329_/B VGND VGND VPWR VPWR _12590_/A sky130_fd_sc_hd__and2_1
XFILLER_114_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12257_ _13716_/A _12257_/B VGND VGND VPWR VPWR _12257_/Y sky130_fd_sc_hd__nor2_1
X_15045_ _15058_/A _15043_/X _15044_/X VGND VGND VPWR VPWR _15045_/X sky130_fd_sc_hd__o21a_1
X_11208_ _13331_/A VGND VGND VPWR VPWR _12215_/A sky130_fd_sc_hd__inv_2
X_12188_ _13716_/A _12257_/B _12187_/Y VGND VGND VPWR VPWR _12188_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11139_ _11136_/Y _12688_/A _10963_/X _11138_/Y VGND VGND VPWR VPWR _11139_/X sky130_fd_sc_hd__o22a_1
X_15947_ _15947_/A _15947_/B VGND VGND VPWR VPWR _15947_/Y sky130_fd_sc_hd__nor2_1
X_15878_ _15878_/A VGND VGND VPWR VPWR _15888_/A sky130_fd_sc_hd__inv_2
XFILLER_63_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14829_ _14742_/X _14772_/A _14771_/X VGND VGND VPWR VPWR _14829_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08350_ _08348_/Y _08349_/A _08348_/A _08349_/Y _08303_/A VGND VGND VPWR VPWR _09221_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08281_ _08281_/A input18/X VGND VGND VPWR VPWR _08282_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ _09856_/B VGND VGND VPWR VPWR _09804_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09735_ _08558_/A _09737_/B _08558_/A _09737_/B VGND VGND VPWR VPWR _09736_/B sky130_fd_sc_hd__a2bb2o_1
X_09666_ _09997_/A _09666_/B VGND VGND VPWR VPWR _09666_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08617_ _08716_/A VGND VGND VPWR VPWR _09456_/A sky130_fd_sc_hd__buf_1
XFILLER_82_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09597_ _09987_/A _09658_/B VGND VGND VPWR VPWR _09597_/Y sky130_fd_sc_hd__nor2_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08690_/A _10118_/B VGND VGND VPWR VPWR _08881_/A sky130_fd_sc_hd__nor2_1
X_08479_ input27/X input11/X VGND VGND VPWR VPWR _08479_/Y sky130_fd_sc_hd__nor2_1
X_11490_ _12393_/A VGND VGND VPWR VPWR _13883_/A sky130_fd_sc_hd__buf_1
X_10510_ _13609_/A VGND VGND VPWR VPWR _11835_/A sky130_fd_sc_hd__inv_2
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10441_ _11028_/A VGND VGND VPWR VPWR _10441_/X sky130_fd_sc_hd__buf_1
XFILLER_7_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13160_ _15252_/A _13113_/B _13113_/Y VGND VGND VPWR VPWR _13160_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10372_ _09117_/A _10371_/X _09117_/A _10371_/X VGND VGND VPWR VPWR _11219_/A sky130_fd_sc_hd__a2bb2o_2
X_12111_ _13196_/A _12061_/B _12061_/Y VGND VGND VPWR VPWR _12111_/Y sky130_fd_sc_hd__o21ai_1
X_13091_ _13011_/X _13090_/X _13011_/X _13090_/X VGND VGND VPWR VPWR _13105_/B sky130_fd_sc_hd__a2bb2o_1
X_12042_ _12042_/A VGND VGND VPWR VPWR _12043_/A sky130_fd_sc_hd__buf_1
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15801_ _15796_/Y _16217_/A _15800_/Y VGND VGND VPWR VPWR _15805_/B sky130_fd_sc_hd__o21ai_1
X_13993_ _13990_/X _13992_/X _13990_/X _13992_/X VGND VGND VPWR VPWR _13995_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15732_ _15544_/A _14920_/B _14920_/Y VGND VGND VPWR VPWR _15732_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12944_ _12944_/A _12944_/B VGND VGND VPWR VPWR _12944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15663_ _15947_/A _15662_/B _14375_/A _14375_/Y _15662_/Y VGND VGND VPWR VPWR _15665_/B
+ sky130_fd_sc_hd__o32a_1
X_12875_ _14677_/A _12942_/B VGND VGND VPWR VPWR _12875_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15594_ _15543_/X _15593_/X _15543_/X _15593_/X VGND VGND VPWR VPWR _15595_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _15345_/A _14660_/B VGND VGND VPWR VPWR _14614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11826_ _11794_/X _11825_/X _11794_/X _11825_/X VGND VGND VPWR VPWR _11837_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14545_/A _14520_/X VGND VGND VPWR VPWR _14545_/X sky130_fd_sc_hd__or2b_1
X_11757_ _11757_/A _11757_/B VGND VGND VPWR VPWR _11757_/X sky130_fd_sc_hd__or2_1
XFILLER_14_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10708_ _11942_/A VGND VGND VPWR VPWR _13068_/A sky130_fd_sc_hd__buf_1
XFILLER_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16215_ _16213_/A _16214_/A _16213_/Y _16214_/Y _16205_/A VGND VGND VPWR VPWR _16253_/A
+ sky130_fd_sc_hd__a221o_1
X_11688_ _11682_/X _11687_/X _11682_/X _11687_/X VGND VGND VPWR VPWR _11688_/Y sky130_fd_sc_hd__o2bb2ai_1
X_14476_ _14471_/X _14475_/X _14471_/X _14475_/X VGND VGND VPWR VPWR _14477_/B sky130_fd_sc_hd__a2bb2o_1
X_13427_ _13423_/Y _13425_/Y _13426_/Y VGND VGND VPWR VPWR _13431_/B sky130_fd_sc_hd__o21ai_1
X_10639_ _10594_/Y _10637_/Y _10638_/Y VGND VGND VPWR VPWR _10640_/A sky130_fd_sc_hd__o21ai_1
XFILLER_127_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16146_ _16119_/A _16119_/B _16119_/Y VGND VGND VPWR VPWR _16148_/A sky130_fd_sc_hd__o21ai_1
X_13358_ _15467_/A _13345_/B _13345_/Y _13357_/X VGND VGND VPWR VPWR _13358_/X sky130_fd_sc_hd__o2bb2a_1
X_16077_ _16038_/A _16038_/B _16038_/Y VGND VGND VPWR VPWR _16077_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12309_ _12309_/A _12309_/B VGND VGND VPWR VPWR _12309_/Y sky130_fd_sc_hd__nand2_1
X_13289_ _13245_/Y _13287_/Y _13288_/Y VGND VGND VPWR VPWR _13290_/A sky130_fd_sc_hd__o21ai_1
X_15028_ _15028_/A _15028_/B VGND VGND VPWR VPWR _15028_/X sky130_fd_sc_hd__or2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput3 wbs_adr_i[10] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_2
X_09520_ _09341_/A _08706_/B _09520_/S VGND VGND VPWR VPWR _09520_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09451_ _09486_/A _09529_/A VGND VGND VPWR VPWR _09451_/Y sky130_fd_sc_hd__nor2_1
X_08402_ _08670_/A VGND VGND VPWR VPWR _08402_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09382_ _10240_/A VGND VGND VPWR VPWR _09383_/B sky130_fd_sc_hd__buf_1
X_08333_ _08333_/A VGND VGND VPWR VPWR _08333_/Y sky130_fd_sc_hd__inv_2
X_08264_ input13/X VGND VGND VPWR VPWR _08346_/B sky130_fd_sc_hd__inv_2
XFILLER_118_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09718_ _09963_/A _10595_/A _09717_/X VGND VGND VPWR VPWR _09720_/B sky130_fd_sc_hd__o21ai_1
X_10990_ _09396_/A _11128_/B _09396_/A _11128_/B VGND VGND VPWR VPWR _10990_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09649_ _09648_/A _09648_/B _09546_/A _09546_/Y _09648_/Y VGND VGND VPWR VPWR _10722_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12660_ _12660_/A VGND VGND VPWR VPWR _12660_/Y sky130_fd_sc_hd__inv_2
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11611_/A VGND VGND VPWR VPWR _11611_/X sky130_fd_sc_hd__buf_1
XFILLER_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14330_ _14388_/A _15958_/A VGND VGND VPWR VPWR _15612_/A sky130_fd_sc_hd__and2_1
X_12591_ _12591_/A VGND VGND VPWR VPWR _12591_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11542_ _11632_/A _11541_/Y _11632_/A _11541_/Y VGND VGND VPWR VPWR _11638_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14261_ _14216_/Y _14259_/Y _14260_/Y VGND VGND VPWR VPWR _14262_/A sky130_fd_sc_hd__o21ai_2
XFILLER_109_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11473_ _09430_/B _09371_/B _09371_/X VGND VGND VPWR VPWR _11474_/B sky130_fd_sc_hd__a21boi_1
X_16000_ _15963_/X _15999_/X _15963_/X _15999_/X VGND VGND VPWR VPWR _16046_/B sky130_fd_sc_hd__a2bb2o_1
X_14192_ _15860_/A _14272_/B VGND VGND VPWR VPWR _14192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13212_ _14841_/A VGND VGND VPWR VPWR _14858_/A sky130_fd_sc_hd__buf_1
X_10424_ _10424_/A _10424_/B VGND VGND VPWR VPWR _10425_/A sky130_fd_sc_hd__or2_1
XFILLER_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13143_ _13124_/X _13142_/Y _13124_/X _13142_/Y VGND VGND VPWR VPWR _13206_/B sky130_fd_sc_hd__a2bb2o_1
X_10355_ _12831_/A _10355_/B VGND VGND VPWR VPWR _10356_/A sky130_fd_sc_hd__nand2_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13074_ _13765_/A VGND VGND VPWR VPWR _15255_/A sky130_fd_sc_hd__buf_1
X_10286_ _13479_/A _10286_/B VGND VGND VPWR VPWR _10289_/A sky130_fd_sc_hd__and2_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12025_ _11971_/X _12024_/Y _11971_/X _12024_/Y VGND VGND VPWR VPWR _12057_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_120_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13976_ _13866_/X _13975_/Y _13876_/Y VGND VGND VPWR VPWR _13998_/A sky130_fd_sc_hd__o21ai_2
X_15715_ _15728_/A _15715_/B VGND VGND VPWR VPWR _16121_/A sky130_fd_sc_hd__or2_1
X_12927_ _12907_/Y _12925_/X _12926_/Y VGND VGND VPWR VPWR _12927_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15646_ _15669_/A _15669_/B VGND VGND VPWR VPWR _15646_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12858_ _12858_/A _12858_/B VGND VGND VPWR VPWR _12858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11809_ _11810_/A _11810_/B VGND VGND VPWR VPWR _11811_/A sky130_fd_sc_hd__and2_1
X_15577_ _14402_/X _15576_/Y _14402_/X _15576_/Y VGND VGND VPWR VPWR _15696_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12789_ _12788_/A _12788_/B _12788_/Y VGND VGND VPWR VPWR _12789_/X sky130_fd_sc_hd__a21o_1
X_14528_ _12001_/Y _14527_/X _12001_/Y _14527_/X VGND VGND VPWR VPWR _14529_/B sky130_fd_sc_hd__o2bb2a_1
X_14459_ _14459_/A _14459_/B VGND VGND VPWR VPWR _14459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16129_ _15987_/X _16128_/X _15987_/X _16128_/X VGND VGND VPWR VPWR _16243_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08951_ _08680_/X _08950_/Y _08680_/X _08950_/Y VGND VGND VPWR VPWR _08951_/Y sky130_fd_sc_hd__a2bb2oi_2
X_08882_ _08689_/X _08881_/Y _08689_/X _08881_/Y VGND VGND VPWR VPWR _08980_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09503_ _09503_/A _09503_/B VGND VGND VPWR VPWR _09503_/Y sky130_fd_sc_hd__nor2_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09434_ _09248_/A _09433_/Y _09426_/Y VGND VGND VPWR VPWR _09436_/B sky130_fd_sc_hd__o21ai_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09365_ _09429_/B _11574_/A VGND VGND VPWR VPWR _09365_/X sky130_fd_sc_hd__or2_1
X_08316_ _08316_/A input20/X VGND VGND VPWR VPWR _08317_/B sky130_fd_sc_hd__nor2_1
X_09296_ _09629_/A _09295_/X _09629_/A _09295_/X VGND VGND VPWR VPWR _09297_/A sky130_fd_sc_hd__a2bb2o_1
X_08247_ input20/X VGND VGND VPWR VPWR _08248_/B sky130_fd_sc_hd__inv_2
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10140_ _10119_/A _10119_/B _10120_/A VGND VGND VPWR VPWR _10143_/A sky130_fd_sc_hd__a21bo_1
XFILLER_102_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10071_ _10071_/A _10071_/B VGND VGND VPWR VPWR _10071_/X sky130_fd_sc_hd__or2_1
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13830_ _13757_/A _13757_/B _13757_/Y VGND VGND VPWR VPWR _13830_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13761_ _13761_/A _13761_/B VGND VGND VPWR VPWR _13761_/X sky130_fd_sc_hd__or2_1
XFILLER_62_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10973_ _10973_/A VGND VGND VPWR VPWR _10973_/Y sky130_fd_sc_hd__inv_2
X_15500_ _15546_/A _15546_/B VGND VGND VPWR VPWR _15500_/X sky130_fd_sc_hd__and2_1
XFILLER_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12712_ _12698_/A _12698_/B _12698_/Y _12711_/X VGND VGND VPWR VPWR _12712_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15431_ _15422_/A _15422_/B _15422_/Y VGND VGND VPWR VPWR _15431_/Y sky130_fd_sc_hd__o21ai_1
X_13692_ _13673_/Y _13690_/X _13691_/Y VGND VGND VPWR VPWR _13692_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12643_ _12643_/A _12643_/B VGND VGND VPWR VPWR _12643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12574_ _12574_/A VGND VGND VPWR VPWR _12574_/Y sky130_fd_sc_hd__inv_2
X_15362_ _15418_/A _15418_/B VGND VGND VPWR VPWR _15438_/A sky130_fd_sc_hd__and2_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14313_ _13440_/A _13440_/B _13440_/Y VGND VGND VPWR VPWR _14313_/X sky130_fd_sc_hd__o21a_1
X_15293_ _15353_/A _15353_/B VGND VGND VPWR VPWR _15357_/A sky130_fd_sc_hd__and2_1
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11525_ rebuffer24/X _11524_/Y _11525_/B1 _11524_/Y VGND VGND VPWR VPWR _11526_/B
+ sky130_fd_sc_hd__a2bb2oi_1
X_14244_ _14244_/A _14244_/B VGND VGND VPWR VPWR _14362_/B sky130_fd_sc_hd__or2_1
XFILLER_109_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11456_ _14120_/A _11377_/B _11377_/Y _12530_/A VGND VGND VPWR VPWR _12522_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14175_ _14128_/X _14174_/Y _14128_/X _14174_/Y VGND VGND VPWR VPWR _14176_/B sky130_fd_sc_hd__a2bb2oi_1
X_11387_ _11391_/A _11387_/B VGND VGND VPWR VPWR _14108_/A sky130_fd_sc_hd__or2_1
X_10407_ _13528_/A _10328_/B _10324_/A _10328_/B VGND VGND VPWR VPWR _10407_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13126_ _13041_/Y _13124_/X _13125_/Y VGND VGND VPWR VPWR _13126_/X sky130_fd_sc_hd__o21a_1
X_10338_ _13530_/A _10338_/B VGND VGND VPWR VPWR _10338_/X sky130_fd_sc_hd__and2_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13057_ _15243_/A _13119_/B VGND VGND VPWR VPWR _13057_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12008_ _12068_/A _12068_/B VGND VGND VPWR VPWR _12008_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10269_ _10234_/Y _10235_/X _10175_/Y _10236_/Y _10472_/A VGND VGND VPWR VPWR _11742_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_78_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13959_ _13897_/Y _13957_/X _13958_/Y VGND VGND VPWR VPWR _13959_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15629_ _14383_/X _15628_/X _14383_/X _15628_/X VGND VGND VPWR VPWR _15673_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09150_ _08512_/X _09146_/X _09150_/S VGND VGND VPWR VPWR _09561_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09081_ _10012_/B _09077_/B _09078_/B VGND VGND VPWR VPWR _09763_/A sky130_fd_sc_hd__a21bo_1
XFILLER_131_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09983_ _09983_/A _09984_/B VGND VGND VPWR VPWR _09983_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08934_ _08934_/A VGND VGND VPWR VPWR _08935_/A sky130_fd_sc_hd__buf_1
X_08865_ _09488_/A _08784_/Y _08786_/Y _08864_/X VGND VGND VPWR VPWR _08865_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08796_ _09209_/A _09453_/B _08713_/X VGND VGND VPWR VPWR _08797_/A sky130_fd_sc_hd__o21ai_1
XFILLER_29_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09417_ _09418_/A _09418_/B VGND VGND VPWR VPWR _09417_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _09525_/A _09348_/B VGND VGND VPWR VPWR _09349_/A sky130_fd_sc_hd__or2_1
XFILLER_21_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11310_ _12266_/A VGND VGND VPWR VPWR _12686_/A sky130_fd_sc_hd__buf_1
X_09279_ _10254_/A VGND VGND VPWR VPWR _09313_/A sky130_fd_sc_hd__buf_1
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12290_ _12290_/A _12358_/B VGND VGND VPWR VPWR _12290_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11241_ _11074_/X _11240_/X _11074_/X _11240_/X VGND VGND VPWR VPWR _11242_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11172_ _11110_/X _11171_/Y _11110_/X _11171_/Y VGND VGND VPWR VPWR _11276_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10123_ _10123_/A _10123_/B VGND VGND VPWR VPWR _10124_/B sky130_fd_sc_hd__or2_1
XFILLER_121_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15980_ _15977_/Y _15979_/X _15977_/Y _15979_/X VGND VGND VPWR VPWR _15982_/B sky130_fd_sc_hd__a2bb2o_1
X_14931_ _14930_/A _14930_/B _14827_/X _14930_/X VGND VGND VPWR VPWR _14931_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10054_ _08930_/A _09505_/Y _08916_/A _09505_/A VGND VGND VPWR VPWR _10055_/B sky130_fd_sc_hd__o22a_1
X_14862_ _14827_/X _14861_/X _14827_/X _14861_/X VGND VGND VPWR VPWR _14928_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13813_ _13813_/A _13767_/X VGND VGND VPWR VPWR _13813_/X sky130_fd_sc_hd__or2b_1
XFILLER_75_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14793_ _14732_/X _14792_/X _14732_/X _14792_/X VGND VGND VPWR VPWR _14794_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13744_ _13761_/A _13761_/B VGND VGND VPWR VPWR _13822_/A sky130_fd_sc_hd__and2_1
XFILLER_44_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10956_ _10956_/A VGND VGND VPWR VPWR _10956_/Y sky130_fd_sc_hd__inv_2
X_16463_ _16357_/A _16463_/D VGND VGND VPWR VPWR _16463_/Q sky130_fd_sc_hd__dfxtp_1
X_10887_ _12051_/A VGND VGND VPWR VPWR _12037_/A sky130_fd_sc_hd__buf_1
X_13675_ _13619_/X _13674_/X _13619_/X _13674_/X VGND VGND VPWR VPWR _13689_/B sky130_fd_sc_hd__a2bb2o_1
X_16394_ _16407_/C _16407_/A VGND VGND VPWR VPWR _16394_/Y sky130_fd_sc_hd__nand2_1
X_12626_ _14208_/A _12624_/X _12625_/X VGND VGND VPWR VPWR _12626_/X sky130_fd_sc_hd__o21a_1
X_15414_ _15414_/A _15414_/B VGND VGND VPWR VPWR _15414_/X sky130_fd_sc_hd__or2_1
XFILLER_31_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15345_ _15345_/A _15345_/B VGND VGND VPWR VPWR _15345_/X sky130_fd_sc_hd__or2_1
XFILLER_12_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12557_ _12557_/A VGND VGND VPWR VPWR _12557_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12488_ _12481_/X _12487_/Y _12481_/X _12487_/Y VGND VGND VPWR VPWR _12488_/X sky130_fd_sc_hd__a2bb2o_1
X_15276_ _14580_/A _15258_/B _15258_/Y _15275_/X VGND VGND VPWR VPWR _15276_/X sky130_fd_sc_hd__a2bb2o_1
X_11508_ _13501_/A _11507_/B _11507_/X _11305_/X VGND VGND VPWR VPWR _11508_/X sky130_fd_sc_hd__o22a_1
X_14227_ _12618_/X _14226_/X _12618_/X _14226_/X VGND VGND VPWR VPWR _14254_/B sky130_fd_sc_hd__a2bb2o_1
X_11439_ _13396_/A VGND VGND VPWR VPWR _15529_/A sky130_fd_sc_hd__buf_1
X_14158_ _14231_/A VGND VGND VPWR VPWR _14207_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13109_ _15258_/A _13109_/B VGND VGND VPWR VPWR _13109_/Y sky130_fd_sc_hd__nand2_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14089_ _14039_/A _14039_/B _13341_/A _14039_/B VGND VGND VPWR VPWR _14089_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08650_ _08650_/A _08650_/B VGND VGND VPWR VPWR _08856_/B sky130_fd_sc_hd__or2_1
XFILLER_94_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08581_ _08580_/X _08428_/X _08580_/X _08428_/X VGND VGND VPWR VPWR _08584_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09202_ _11411_/B VGND VGND VPWR VPWR _11249_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09133_ _09426_/A _09136_/B VGND VGND VPWR VPWR _09133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09064_ _09064_/A VGND VGND VPWR VPWR _09064_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09966_ _10083_/A VGND VGND VPWR VPWR _09966_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09897_/A _09855_/X VGND VGND VPWR VPWR _09898_/B sky130_fd_sc_hd__or2b_1
X_08917_ _08917_/A VGND VGND VPWR VPWR _08922_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _09503_/B _08722_/X _08847_/A _08722_/X VGND VGND VPWR VPWR _08935_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_72_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08779_ _09452_/A VGND VGND VPWR VPWR _09488_/A sky130_fd_sc_hd__buf_1
X_11790_ _10426_/B _11789_/Y _10426_/B _11789_/Y VGND VGND VPWR VPWR _11791_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10810_ _10807_/Y _12692_/A _10672_/X _10809_/Y VGND VGND VPWR VPWR _10810_/X sky130_fd_sc_hd__o22a_1
XFILLER_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10741_ _10741_/A VGND VGND VPWR VPWR _10741_/Y sky130_fd_sc_hd__inv_2
X_13460_ _15171_/A VGND VGND VPWR VPWR _15425_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12411_ _13495_/A VGND VGND VPWR VPWR _13458_/A sky130_fd_sc_hd__buf_1
XFILLER_43_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10672_ _10669_/Y _12694_/A _10553_/X _10671_/Y VGND VGND VPWR VPWR _10672_/X sky130_fd_sc_hd__o22a_1
X_13391_ _13391_/A _13363_/X VGND VGND VPWR VPWR _13391_/X sky130_fd_sc_hd__or2b_1
X_12342_ _12218_/A _12218_/B _12218_/Y VGND VGND VPWR VPWR _12342_/Y sky130_fd_sc_hd__o21ai_1
X_15130_ _15092_/X _15129_/Y _15092_/X _15129_/Y VGND VGND VPWR VPWR _15131_/B sky130_fd_sc_hd__a2bb2o_1
X_15061_ _15061_/A _15042_/X VGND VGND VPWR VPWR _15061_/X sky130_fd_sc_hd__or2b_1
X_12273_ _12273_/A _12273_/B VGND VGND VPWR VPWR _12273_/X sky130_fd_sc_hd__or2_1
XFILLER_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11224_ _12221_/A _11224_/B VGND VGND VPWR VPWR _11224_/Y sky130_fd_sc_hd__nand2_1
X_14012_ _14012_/A _14062_/B VGND VGND VPWR VPWR _14129_/A sky130_fd_sc_hd__and2_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11155_ _11155_/A _11155_/B VGND VGND VPWR VPWR _11155_/Y sky130_fd_sc_hd__nand2_1
X_15963_ _16002_/A _15961_/X _15962_/X VGND VGND VPWR VPWR _15963_/X sky130_fd_sc_hd__o21a_1
X_11086_ _11216_/A _11084_/X _11085_/X VGND VGND VPWR VPWR _11086_/X sky130_fd_sc_hd__o21a_1
X_10106_ _10177_/A _10177_/B VGND VGND VPWR VPWR _10106_/Y sky130_fd_sc_hd__nand2_1
X_14914_ _14914_/A _14914_/B VGND VGND VPWR VPWR _14914_/Y sky130_fd_sc_hd__nand2_1
X_10037_ _10087_/A _10087_/B VGND VGND VPWR VPWR _10037_/X sky130_fd_sc_hd__and2_1
X_15894_ _15894_/A _15894_/B VGND VGND VPWR VPWR _15894_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14845_ _14944_/A _14944_/B _14844_/Y VGND VGND VPWR VPWR _14845_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14776_ _14776_/A _14741_/X VGND VGND VPWR VPWR _14776_/X sky130_fd_sc_hd__or2b_1
X_11988_ _11988_/A VGND VGND VPWR VPWR _12075_/A sky130_fd_sc_hd__inv_2
XFILLER_44_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13727_ _13727_/A _13701_/X VGND VGND VPWR VPWR _13727_/X sky130_fd_sc_hd__or2b_1
XFILLER_44_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10939_ _10939_/A VGND VGND VPWR VPWR _10939_/Y sky130_fd_sc_hd__inv_2
X_16446_ _16471_/Q VGND VGND VPWR VPWR _16446_/Y sky130_fd_sc_hd__inv_2
X_13658_ _13701_/A _13701_/B VGND VGND VPWR VPWR _13727_/A sky130_fd_sc_hd__and2_1
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16377_ _08230_/A _16460_/Q _08233_/A _16397_/A _16343_/A VGND VGND VPWR VPWR _16460_/D
+ sky130_fd_sc_hd__o221a_2
X_12609_ _12609_/A VGND VGND VPWR VPWR _12610_/A sky130_fd_sc_hd__buf_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13589_ _13580_/X _13588_/Y _13580_/X _13588_/Y VGND VGND VPWR VPWR _13638_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15328_ _11064_/B _15327_/X _11064_/B _15327_/X VGND VGND VPWR VPWR _15329_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15259_ _15205_/A _15205_/B _15205_/Y VGND VGND VPWR VPWR _15259_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09820_ _09820_/A _09820_/B VGND VGND VPWR VPWR _09821_/B sky130_fd_sc_hd__or2_1
XFILLER_101_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09751_ _09745_/A _09745_/B _09791_/A VGND VGND VPWR VPWR _10087_/A sky130_fd_sc_hd__a21bo_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ _08703_/A _09146_/A VGND VGND VPWR VPWR _09341_/A sky130_fd_sc_hd__nor2_1
XFILLER_94_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09682_ _08657_/A _09684_/B _08657_/A _09684_/B VGND VGND VPWR VPWR _09683_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08633_ _08632_/X _08408_/Y _08632_/X _08408_/Y VGND VGND VPWR VPWR _08635_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08564_ _09453_/B VGND VGND VPWR VPWR _09555_/A sky130_fd_sc_hd__buf_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08495_ _08242_/A _08306_/B _08469_/Y _08501_/A VGND VGND VPWR VPWR _08699_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09116_ _09547_/B _09032_/B _09033_/B VGND VGND VPWR VPWR _09117_/A sky130_fd_sc_hd__a21bo_1
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09047_ _09047_/A VGND VGND VPWR VPWR _09047_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09949_ _09949_/A VGND VGND VPWR VPWR _11770_/A sky130_fd_sc_hd__buf_1
XFILLER_85_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12960_ _12943_/X _12959_/Y _12943_/X _12959_/Y VGND VGND VPWR VPWR _13032_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12891_ _14469_/A _12934_/B VGND VGND VPWR VPWR _12891_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11911_ _13552_/A _11911_/B VGND VGND VPWR VPWR _11911_/X sky130_fd_sc_hd__and2_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _15337_/A _14652_/B VGND VGND VPWR VPWR _14630_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11842_ _11821_/Y _11840_/X _11841_/Y VGND VGND VPWR VPWR _11842_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14561_/A _14512_/X VGND VGND VPWR VPWR _14561_/X sky130_fd_sc_hd__or2b_1
XFILLER_54_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16324_/A _16258_/B _16258_/Y VGND VGND VPWR VPWR _16300_/Y sky130_fd_sc_hd__o21ai_1
X_11773_ _12767_/A _11772_/B _11772_/Y VGND VGND VPWR VPWR _11773_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13512_ _10692_/X _13487_/X _10692_/X _13487_/X VGND VGND VPWR VPWR _13513_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _15202_/A _14516_/B VGND VGND VPWR VPWR _14553_/A sky130_fd_sc_hd__and2_1
X_10724_ _10722_/A _10723_/A _10722_/Y _10723_/Y _09672_/A VGND VGND VPWR VPWR _11970_/A
+ sky130_fd_sc_hd__a221o_2
X_16231_ _16251_/A _16231_/B VGND VGND VPWR VPWR _16231_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13443_ _13387_/Y _13441_/X _13442_/Y VGND VGND VPWR VPWR _13443_/X sky130_fd_sc_hd__o21a_1
X_10655_ _10653_/Y _10654_/Y _10654_/B _09906_/X _10792_/A VGND VGND VPWR VPWR _12936_/A
+ sky130_fd_sc_hd__o221a_2
X_16162_ _16268_/A _16334_/A VGND VGND VPWR VPWR _16162_/Y sky130_fd_sc_hd__nor2_1
X_13374_ _13310_/X _13373_/X _13310_/X _13373_/X VGND VGND VPWR VPWR _13450_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12325_ _15512_/A _12322_/B _12322_/X _12600_/A VGND VGND VPWR VPWR _12329_/B sky130_fd_sc_hd__o22a_1
X_15113_ _15113_/A _15113_/B VGND VGND VPWR VPWR _15113_/Y sky130_fd_sc_hd__nand2_1
X_10586_ _11843_/A _10533_/B _10533_/Y VGND VGND VPWR VPWR _10586_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16093_ _16031_/X _16092_/Y _16031_/X _16092_/Y VGND VGND VPWR VPWR _16213_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12256_ _12254_/Y _12255_/Y _12190_/Y VGND VGND VPWR VPWR _12363_/A sky130_fd_sc_hd__o21ai_1
X_15044_ _15044_/A _15044_/B VGND VGND VPWR VPWR _15044_/X sky130_fd_sc_hd__or2_1
XFILLER_5_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11207_ _11207_/A _11219_/B VGND VGND VPWR VPWR _13331_/A sky130_fd_sc_hd__or2_1
X_12187_ _12187_/A _12257_/B VGND VGND VPWR VPWR _12187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11138_ _11138_/A _12087_/A VGND VGND VPWR VPWR _11138_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15946_ _14371_/X _14373_/Y _15839_/B _14375_/A _14370_/A VGND VGND VPWR VPWR _15947_/B
+ sky130_fd_sc_hd__o221a_1
X_11069_ _12135_/A VGND VGND VPWR VPWR _14430_/A sky130_fd_sc_hd__buf_1
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15877_ _15890_/A _15890_/B VGND VGND VPWR VPWR _15877_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14828_ _15437_/A VGND VGND VPWR VPWR _14930_/A sky130_fd_sc_hd__buf_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14759_ _14750_/X _14758_/X _14750_/X _14758_/X VGND VGND VPWR VPWR _14761_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08280_ input2/X VGND VGND VPWR VPWR _08358_/A sky130_fd_sc_hd__inv_2
XFILLER_32_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16429_ _16447_/A _16429_/B VGND VGND VPWR VPWR _16429_/X sky130_fd_sc_hd__or2_1
XFILLER_20_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09803_ _09803_/A _09803_/B VGND VGND VPWR VPWR _09856_/B sky130_fd_sc_hd__or2_1
XFILLER_101_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09734_ _09734_/A _09734_/B VGND VGND VPWR VPWR _09737_/B sky130_fd_sc_hd__or2_1
XFILLER_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09665_ _09579_/Y _09663_/X _09664_/Y VGND VGND VPWR VPWR _09665_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08616_ _09221_/A VGND VGND VPWR VPWR _08716_/A sky130_fd_sc_hd__inv_2
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09596_ _09554_/X _09595_/Y _09554_/X _09595_/Y VGND VGND VPWR VPWR _09658_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08547_ _08546_/A _08446_/Y _08546_/Y _08446_/A VGND VGND VPWR VPWR _10118_/B sky130_fd_sc_hd__o22a_1
X_08478_ input28/X input12/X VGND VGND VPWR VPWR _08478_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10440_ _10438_/A _10439_/A _10438_/Y _10439_/Y _09393_/A VGND VGND VPWR VPWR _11028_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10371_ _09415_/A _09118_/B _09118_/Y VGND VGND VPWR VPWR _10371_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12110_ _13902_/A _12151_/B VGND VGND VPWR VPWR _12207_/A sky130_fd_sc_hd__and2_1
X_13090_ _13090_/A _13013_/X VGND VGND VPWR VPWR _13090_/X sky130_fd_sc_hd__or2b_1
XFILLER_123_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12041_ _12041_/A _12041_/B VGND VGND VPWR VPWR _12042_/A sky130_fd_sc_hd__or2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15800_ _16099_/A _15800_/B VGND VGND VPWR VPWR _15800_/Y sky130_fd_sc_hd__nand2_1
X_13992_ _13861_/X _13991_/Y _13886_/Y VGND VGND VPWR VPWR _13992_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15731_ _16114_/A _15815_/B VGND VGND VPWR VPWR _15731_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12943_ _12875_/Y _12941_/X _12942_/Y VGND VGND VPWR VPWR _12943_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15662_ _15947_/A _15662_/B VGND VGND VPWR VPWR _15662_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12874_ _12855_/X _12873_/Y _12855_/X _12873_/Y VGND VGND VPWR VPWR _12942_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15593_ _15503_/X _15593_/B VGND VGND VPWR VPWR _15593_/X sky130_fd_sc_hd__and2b_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _14587_/X _14612_/Y _14587_/X _14612_/Y VGND VGND VPWR VPWR _14660_/B sky130_fd_sc_hd__a2bb2o_1
X_11825_ _11780_/A _11780_/B _11780_/A _11780_/B VGND VGND VPWR VPWR _11825_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _15252_/A VGND VGND VPWR VPWR _14584_/A sky130_fd_sc_hd__buf_1
X_11756_ _11798_/A VGND VGND VPWR VPWR _12769_/A sky130_fd_sc_hd__buf_1
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _14474_/A _14474_/B _14474_/Y VGND VGND VPWR VPWR _14475_/X sky130_fd_sc_hd__a21o_1
X_10707_ _10930_/A _10707_/B VGND VGND VPWR VPWR _11942_/A sky130_fd_sc_hd__or2_2
XFILLER_14_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16214_ _16214_/A VGND VGND VPWR VPWR _16214_/Y sky130_fd_sc_hd__inv_2
X_13426_ _14101_/A _13426_/B VGND VGND VPWR VPWR _13426_/Y sky130_fd_sc_hd__nand2_1
X_11687_ _11684_/X _11686_/X _11684_/X _11686_/X VGND VGND VPWR VPWR _11687_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_127_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10638_ _11901_/A _10638_/B VGND VGND VPWR VPWR _10638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16145_ _16273_/A _16272_/A VGND VGND VPWR VPWR _16145_/Y sky130_fd_sc_hd__nor2_1
X_13357_ _15470_/A _13349_/B _13349_/Y _13356_/Y VGND VGND VPWR VPWR _13357_/X sky130_fd_sc_hd__o2bb2a_1
X_10569_ _10569_/A _10569_/B VGND VGND VPWR VPWR _10569_/Y sky130_fd_sc_hd__nand2_1
X_16076_ _16108_/A _16108_/B VGND VGND VPWR VPWR _16076_/X sky130_fd_sc_hd__and2_1
XFILLER_115_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12308_ _12244_/X _12307_/Y _12244_/X _12307_/Y VGND VGND VPWR VPWR _12309_/B sky130_fd_sc_hd__a2bb2o_1
X_13288_ _14733_/A _13288_/B VGND VGND VPWR VPWR _13288_/Y sky130_fd_sc_hd__nand2_1
X_12239_ _13341_/A _12227_/B _12227_/Y _12238_/X VGND VGND VPWR VPWR _12239_/X sky130_fd_sc_hd__a2bb2o_1
X_15027_ _12829_/A _12829_/B _10426_/A _12829_/Y VGND VGND VPWR VPWR _15027_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 wbs_adr_i[11] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_4
X_15929_ _15895_/X _15928_/Y _15895_/X _15928_/Y VGND VGND VPWR VPWR _15958_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09450_ _09484_/A _09527_/A VGND VGND VPWR VPWR _09450_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08401_ _08401_/A _09677_/B VGND VGND VPWR VPWR _08670_/A sky130_fd_sc_hd__or2_1
XFILLER_101_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09381_ _09335_/X _08883_/Y _09335_/X _08883_/Y VGND VGND VPWR VPWR _10240_/A sky130_fd_sc_hd__o2bb2a_1
X_08332_ _08332_/A _08332_/B VGND VGND VPWR VPWR _08333_/A sky130_fd_sc_hd__or2_1
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08263_ _08263_/A input14/X VGND VGND VPWR VPWR _08342_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09717_ _09717_/A _09717_/B VGND VGND VPWR VPWR _09717_/X sky130_fd_sc_hd__or2_1
XFILLER_55_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09648_ _09648_/A _09648_/B VGND VGND VPWR VPWR _09648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09995_/A _09664_/B VGND VGND VPWR VPWR _09579_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12590_ _12590_/A _12329_/X VGND VGND VPWR VPWR _12591_/A sky130_fd_sc_hd__or2b_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11609_/A _12423_/B _11609_/Y VGND VGND VPWR VPWR _11611_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11541_ _12440_/A _11631_/B _11540_/Y VGND VGND VPWR VPWR _11541_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14260_ _15872_/A _14260_/B VGND VGND VPWR VPWR _14260_/Y sky130_fd_sc_hd__nand2_1
X_11472_ _11351_/A _11267_/X _11350_/X VGND VGND VPWR VPWR _11472_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14191_ _12630_/X _14190_/X _12630_/X _14190_/X VGND VGND VPWR VPWR _14272_/B sky130_fd_sc_hd__a2bb2o_1
X_13211_ _15107_/A VGND VGND VPWR VPWR _14841_/A sky130_fd_sc_hd__inv_2
X_10423_ _10423_/A VGND VGND VPWR VPWR _10424_/B sky130_fd_sc_hd__inv_2
XFILLER_124_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13142_ _14953_/A _13125_/B _13125_/Y VGND VGND VPWR VPWR _13142_/Y sky130_fd_sc_hd__o21ai_1
X_10354_ _10424_/A _10421_/B VGND VGND VPWR VPWR _10354_/X sky130_fd_sc_hd__or2_1
XFILLER_3_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13073_ _13073_/A VGND VGND VPWR VPWR _13765_/A sky130_fd_sc_hd__inv_2
X_10285_ _10282_/A _10281_/A _10350_/A _10284_/Y VGND VGND VPWR VPWR _10286_/B sky130_fd_sc_hd__o22a_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12024_ _13073_/A _11972_/B _11972_/Y VGND VGND VPWR VPWR _12024_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13975_ _13975_/A _13975_/B VGND VGND VPWR VPWR _13975_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15714_ _14925_/X _15713_/X _14925_/X _15713_/X VGND VGND VPWR VPWR _15715_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_73_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12926_ _12926_/A _12926_/B VGND VGND VPWR VPWR _12926_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15645_ _14379_/X _15644_/X _14379_/X _15644_/X VGND VGND VPWR VPWR _15669_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12857_ _12798_/Y _12855_/X _12856_/Y VGND VGND VPWR VPWR _12857_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11808_ _10467_/A _11807_/A _10467_/Y _11854_/B VGND VGND VPWR VPWR _11810_/B sky130_fd_sc_hd__o22a_1
X_15576_ _15972_/A _14403_/B _14403_/Y VGND VGND VPWR VPWR _15576_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _12788_/A _12788_/B VGND VGND VPWR VPWR _12788_/Y sky130_fd_sc_hd__nor2_1
X_11739_ _11777_/B VGND VGND VPWR VPWR _11739_/Y sky130_fd_sc_hd__inv_2
X_14527_ _15040_/A _11986_/Y _11928_/Y _14472_/X VGND VGND VPWR VPWR _14527_/X sky130_fd_sc_hd__o22a_1
X_14458_ _13610_/Y _13616_/A _13617_/Y VGND VGND VPWR VPWR _14458_/Y sky130_fd_sc_hd__o21ai_1
X_14389_ _15612_/A _14387_/X _14388_/X VGND VGND VPWR VPWR _14389_/X sky130_fd_sc_hd__o21a_1
X_13409_ _15470_/A _13349_/B _13349_/Y VGND VGND VPWR VPWR _13409_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16128_ _16126_/Y _16127_/X _16126_/Y _16127_/X VGND VGND VPWR VPWR _16128_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_115_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16059_ _16059_/A _16055_/X VGND VGND VPWR VPWR _16059_/X sky130_fd_sc_hd__or2b_1
X_08950_ _09539_/A _08647_/A _08648_/X VGND VGND VPWR VPWR _08950_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08881_ _08881_/A _08881_/B VGND VGND VPWR VPWR _08881_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09502_ _09502_/A _09502_/B VGND VGND VPWR VPWR _09502_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09433_ _09766_/A _09433_/B VGND VGND VPWR VPWR _09433_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _08753_/Y _09338_/Y _08753_/Y _09338_/Y VGND VGND VPWR VPWR _11574_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_52_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08315_ _08313_/Y _08314_/A _08313_/A _08314_/Y _08304_/X VGND VGND VPWR VPWR _08532_/B
+ sky130_fd_sc_hd__o221a_1
X_09295_ _09502_/A _09006_/Y _09540_/A _09231_/Y VGND VGND VPWR VPWR _09295_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08246_ input4/X VGND VGND VPWR VPWR _08316_/A sky130_fd_sc_hd__inv_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10070_ _10022_/X _10069_/Y _10022_/X _10069_/Y VGND VGND VPWR VPWR _10071_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13760_ _13826_/A _13758_/X _13759_/X VGND VGND VPWR VPWR _13760_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10972_ _10972_/A VGND VGND VPWR VPWR _10972_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13691_ _14493_/A _13691_/B VGND VGND VPWR VPWR _13691_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12711_ _12700_/A _12700_/B _12700_/Y _12710_/X VGND VGND VPWR VPWR _12711_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12642_ _11671_/X _12642_/B VGND VGND VPWR VPWR _12643_/B sky130_fd_sc_hd__and2b_1
X_15430_ _14971_/A _15167_/B _15167_/Y _15169_/Y VGND VGND VPWR VPWR _15430_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12573_ _12623_/A _12623_/B VGND VGND VPWR VPWR _14214_/A sky130_fd_sc_hd__and2_1
X_15361_ _15350_/X _15360_/X _15350_/X _15360_/X VGND VGND VPWR VPWR _15418_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14312_ _15964_/A _14394_/B VGND VGND VPWR VPWR _15590_/A sky130_fd_sc_hd__and2_1
X_15292_ _15283_/X _15291_/Y _15283_/X _15291_/Y VGND VGND VPWR VPWR _15353_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11524_ _10238_/B _10139_/B _10139_/Y VGND VGND VPWR VPWR _11524_/Y sky130_fd_sc_hd__a21oi_1
X_14243_ _14243_/A _14243_/B VGND VGND VPWR VPWR _14372_/B sky130_fd_sc_hd__nor2_1
X_11455_ _14114_/A _11384_/B _11384_/Y _12538_/A VGND VGND VPWR VPWR _12530_/A sky130_fd_sc_hd__a2bb2o_1
X_10406_ _11780_/A VGND VGND VPWR VPWR _13568_/A sky130_fd_sc_hd__buf_1
XFILLER_109_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14174_ _13444_/A _14133_/A _14131_/Y VGND VGND VPWR VPWR _14174_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11386_ _08971_/X _11385_/X _08971_/X _11385_/X VGND VGND VPWR VPWR _11387_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13125_ _15234_/A _13125_/B VGND VGND VPWR VPWR _13125_/Y sky130_fd_sc_hd__nand2_1
X_10337_ _10291_/B _10336_/Y _10291_/B _10336_/Y VGND VGND VPWR VPWR _10338_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13056_ _13027_/X _13055_/X _13027_/X _13055_/X VGND VGND VPWR VPWR _13119_/B sky130_fd_sc_hd__a2bb2o_1
X_10268_ _10268_/A VGND VGND VPWR VPWR _10472_/A sky130_fd_sc_hd__clkbuf_2
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12007_ _11982_/X _12006_/Y _11982_/X _12006_/Y VGND VGND VPWR VPWR _12068_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10199_ _10196_/X _10198_/X _10196_/X _10198_/X VGND VGND VPWR VPWR _10346_/B sky130_fd_sc_hd__o2bb2a_4
XFILLER_66_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13958_ _15416_/A _13958_/B VGND VGND VPWR VPWR _13958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12909_ _15084_/A _12838_/B _12838_/Y VGND VGND VPWR VPWR _12909_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13889_ _15420_/A _13962_/B VGND VGND VPWR VPWR _13889_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15628_ _15628_/A _14384_/X VGND VGND VPWR VPWR _15628_/X sky130_fd_sc_hd__or2b_1
XFILLER_15_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15559_ _15430_/X _15558_/X _15430_/X _15558_/X VGND VGND VPWR VPWR _15559_/X sky130_fd_sc_hd__a2bb2o_1
X_09080_ _09760_/A VGND VGND VPWR VPWR _09432_/A sky130_fd_sc_hd__buf_1
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09982_ _09700_/Y _09980_/Y _09981_/Y VGND VGND VPWR VPWR _09984_/B sky130_fd_sc_hd__o21ai_1
XFILLER_130_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08933_ _10228_/B _08932_/B _08931_/Y _08932_/Y VGND VGND VPWR VPWR _08942_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08864_ _09490_/A _08792_/Y _08793_/Y _08863_/X VGND VGND VPWR VPWR _08864_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08795_ _09492_/A VGND VGND VPWR VPWR _08795_/X sky130_fd_sc_hd__buf_1
XFILLER_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09416_ _09946_/A _09414_/Y _09415_/Y VGND VGND VPWR VPWR _09418_/B sky130_fd_sc_hd__o21ai_1
X_09347_ _09347_/A VGND VGND VPWR VPWR _09347_/Y sky130_fd_sc_hd__inv_2
X_09278_ _09257_/X _08910_/Y _09257_/X _08910_/Y VGND VGND VPWR VPWR _10254_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08229_ _08229_/A VGND VGND VPWR VPWR _08230_/A sky130_fd_sc_hd__buf_1
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11240_ _11240_/A _11076_/X VGND VGND VPWR VPWR _11240_/X sky130_fd_sc_hd__or2b_1
XFILLER_106_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11171_ _13048_/A _11170_/B _11170_/Y VGND VGND VPWR VPWR _11171_/Y sky130_fd_sc_hd__o21ai_1
X_10122_ _10237_/B VGND VGND VPWR VPWR _10122_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14930_ _14930_/A _14930_/B VGND VGND VPWR VPWR _14930_/X sky130_fd_sc_hd__and2_1
XFILLER_88_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10053_ _09066_/A _09681_/A _09401_/Y _08931_/A VGND VGND VPWR VPWR _10055_/A sky130_fd_sc_hd__o22a_1
X_14861_ _14930_/A _14930_/B _14930_/A _14930_/B VGND VGND VPWR VPWR _14861_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13812_ _14615_/A _13852_/B VGND VGND VPWR VPWR _13812_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14792_ _14792_/A _14733_/X VGND VGND VPWR VPWR _14792_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13743_ _13690_/X _13742_/Y _13690_/X _13742_/Y VGND VGND VPWR VPWR _13761_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10955_ _09990_/A _09990_/B _09990_/Y VGND VGND VPWR VPWR _10956_/A sky130_fd_sc_hd__o21ai_1
X_16462_ _16357_/A _16462_/D VGND VGND VPWR VPWR _16462_/Q sky130_fd_sc_hd__dfxtp_1
X_13674_ _15140_/A _13606_/B _13606_/Y VGND VGND VPWR VPWR _13674_/X sky130_fd_sc_hd__a21o_1
X_10886_ _10402_/A _10885_/Y _10402_/Y _10885_/A _09445_/A VGND VGND VPWR VPWR _12051_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16393_ _16402_/A VGND VGND VPWR VPWR _16393_/Y sky130_fd_sc_hd__inv_2
X_12625_ _12625_/A _12625_/B VGND VGND VPWR VPWR _12625_/X sky130_fd_sc_hd__or2_1
X_15413_ _15447_/A _15411_/X _15412_/X VGND VGND VPWR VPWR _15413_/X sky130_fd_sc_hd__o21a_1
X_12556_ _14914_/A _11446_/B _11446_/Y VGND VGND VPWR VPWR _12557_/A sky130_fd_sc_hd__o21ai_1
X_15344_ _15372_/A _15342_/X _15343_/X VGND VGND VPWR VPWR _15344_/X sky130_fd_sc_hd__o21a_1
X_11507_ _13501_/A _11507_/B VGND VGND VPWR VPWR _11507_/X sky130_fd_sc_hd__and2_1
XFILLER_8_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12487_ _12484_/Y _12485_/Y _12486_/Y VGND VGND VPWR VPWR _12487_/Y sky130_fd_sc_hd__o21ai_1
X_15275_ _14578_/A _15261_/B _15261_/Y _15274_/X VGND VGND VPWR VPWR _15275_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14226_ _14226_/A _12619_/X VGND VGND VPWR VPWR _14226_/X sky130_fd_sc_hd__or2b_1
X_11438_ _11254_/X _11437_/Y _11254_/X _11437_/Y VGND VGND VPWR VPWR _12564_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14157_ _14245_/A VGND VGND VPWR VPWR _14231_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11369_ _11259_/X _11368_/Y _11259_/X _11368_/Y VGND VGND VPWR VPWR _11370_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13108_ _13087_/Y _13106_/X _13107_/Y VGND VGND VPWR VPWR _13108_/X sky130_fd_sc_hd__o21a_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14088_ _14091_/A _14091_/B VGND VGND VPWR VPWR _14088_/X sky130_fd_sc_hd__and2_1
XFILLER_79_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _13039_/A _13034_/X VGND VGND VPWR VPWR _13039_/X sky130_fd_sc_hd__or2b_1
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08580_ _09324_/A _09209_/B _10013_/A _08579_/Y VGND VGND VPWR VPWR _08580_/X sky130_fd_sc_hd__o22a_1
XFILLER_93_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09201_ _09193_/Y _09200_/X _09193_/Y _09200_/X VGND VGND VPWR VPWR _11411_/B sky130_fd_sc_hd__a2bb2o_4
X_09132_ _09128_/Y _09130_/Y _09131_/Y VGND VGND VPWR VPWR _09136_/B sky130_fd_sc_hd__o21ai_2
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09063_ _08839_/A _09042_/X _08839_/A _09042_/X VGND VGND VPWR VPWR _09070_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09965_ _09995_/A _09995_/B VGND VGND VPWR VPWR _09965_/X sky130_fd_sc_hd__and2_1
XFILLER_97_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _09882_/A _09882_/B _09883_/B VGND VGND VPWR VPWR _09898_/A sky130_fd_sc_hd__a21bo_1
X_08916_ _08916_/A _09817_/B VGND VGND VPWR VPWR _08917_/A sky130_fd_sc_hd__or2_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _08847_/A VGND VGND VPWR VPWR _09503_/B sky130_fd_sc_hd__buf_1
XFILLER_18_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08778_ _08778_/A _08778_/B VGND VGND VPWR VPWR _08778_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10740_ _10740_/A VGND VGND VPWR VPWR _10740_/Y sky130_fd_sc_hd__inv_2
X_10671_ _10671_/A _11859_/A VGND VGND VPWR VPWR _10671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12410_ _12410_/A VGND VGND VPWR VPWR _13495_/A sky130_fd_sc_hd__buf_1
XFILLER_9_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13390_ _14120_/A _13440_/B VGND VGND VPWR VPWR _13390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12341_ _12344_/A _12344_/B VGND VGND VPWR VPWR _12341_/Y sky130_fd_sc_hd__nor2_1
X_15060_ _15060_/A _15060_/B VGND VGND VPWR VPWR _15060_/Y sky130_fd_sc_hd__nand2_1
X_12272_ _12273_/A _12273_/B VGND VGND VPWR VPWR _12274_/A sky130_fd_sc_hd__and2_1
XFILLER_122_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14011_ _13957_/X _14010_/Y _13957_/X _14010_/Y VGND VGND VPWR VPWR _14062_/B sky130_fd_sc_hd__a2bb2o_1
X_11223_ _11082_/X _11222_/X _11082_/X _11222_/X VGND VGND VPWR VPWR _11224_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11154_ _09383_/B _10240_/B _10240_/X VGND VGND VPWR VPWR _11155_/B sky130_fd_sc_hd__a21boi_1
X_15962_ _15962_/A _15962_/B VGND VGND VPWR VPWR _15962_/X sky130_fd_sc_hd__or2_1
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11085_ _13914_/A _11085_/B VGND VGND VPWR VPWR _11085_/X sky130_fd_sc_hd__or2_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10105_ _08671_/A _08667_/A _09627_/A _08667_/Y VGND VGND VPWR VPWR _10177_/B sky130_fd_sc_hd__o22a_1
X_14913_ _14892_/Y _14911_/X _14912_/Y VGND VGND VPWR VPWR _14913_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10036_ _10029_/X _10035_/Y _10029_/X _10035_/Y VGND VGND VPWR VPWR _10087_/B sky130_fd_sc_hd__a2bb2o_1
X_15893_ _15874_/Y _15891_/X _15892_/Y VGND VGND VPWR VPWR _15893_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14844_ _14944_/A _14944_/B VGND VGND VPWR VPWR _14844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14775_ _15443_/A VGND VGND VPWR VPWR _14778_/A sky130_fd_sc_hd__buf_1
XFILLER_91_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11987_ _11985_/A _11985_/B _11985_/X _11986_/Y VGND VGND VPWR VPWR _12075_/B sky130_fd_sc_hd__a22o_1
XFILLER_17_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13726_ _13773_/A _13773_/B VGND VGND VPWR VPWR _13804_/A sky130_fd_sc_hd__and2_1
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10938_ _09779_/A _09779_/B _09779_/Y VGND VGND VPWR VPWR _10939_/A sky130_fd_sc_hd__o21ai_1
X_16445_ _16445_/A _16445_/B VGND VGND VPWR VPWR _16445_/X sky130_fd_sc_hd__and2_1
XFILLER_71_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13657_ _13640_/A _13656_/Y _13640_/A _13656_/Y VGND VGND VPWR VPWR _13701_/B sky130_fd_sc_hd__a2bb2o_1
X_10869_ _10869_/A VGND VGND VPWR VPWR _10869_/Y sky130_fd_sc_hd__inv_2
X_16376_ _16319_/X _16375_/Y _16319_/X _16375_/Y VGND VGND VPWR VPWR _16397_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12608_ _14244_/A _12607_/B _12607_/Y _11705_/A VGND VGND VPWR VPWR _14235_/A sky130_fd_sc_hd__o211a_1
X_13588_ _13548_/A _13548_/B _13549_/A VGND VGND VPWR VPWR _13588_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12539_ _12538_/A _12538_/B _12538_/Y _11707_/A VGND VGND VPWR VPWR _12629_/A sky130_fd_sc_hd__o211a_1
X_15327_ _14568_/A _15270_/B _14568_/A _15270_/B VGND VGND VPWR VPWR _15327_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15258_ _15258_/A _15258_/B VGND VGND VPWR VPWR _15258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14209_ _12624_/X _14208_/X _12624_/X _14208_/X VGND VGND VPWR VPWR _14263_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15189_ _15154_/X _15188_/Y _15154_/X _15188_/Y VGND VGND VPWR VPWR _15190_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09750_ _09750_/A _09750_/B VGND VGND VPWR VPWR _09750_/Y sky130_fd_sc_hd__nor2_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ _08701_/A _08701_/B VGND VGND VPWR VPWR _08703_/A sky130_fd_sc_hd__or2_2
X_09681_ _09681_/A _09681_/B VGND VGND VPWR VPWR _09684_/B sky130_fd_sc_hd__or2_1
XFILLER_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08632_ _09252_/A _09225_/B _10017_/A _08631_/Y VGND VGND VPWR VPWR _08632_/X sky130_fd_sc_hd__o22a_1
XFILLER_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08563_ _08589_/A _08563_/B VGND VGND VPWR VPWR _09453_/B sky130_fd_sc_hd__or2_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08494_ _08311_/A _08245_/B _08470_/Y _08516_/A VGND VGND VPWR VPWR _08501_/A sky130_fd_sc_hd__o22a_1
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09115_ _09415_/A _09118_/B VGND VGND VPWR VPWR _09115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09046_ _08715_/A _08715_/B _08715_/X _09045_/X VGND VGND VPWR VPWR _09047_/A sky130_fd_sc_hd__a22o_1
XFILLER_116_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09948_ _09946_/A _09947_/A _09946_/Y _09947_/Y _09392_/A VGND VGND VPWR VPWR _09949_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09879_ _09867_/X _08789_/Y _09867_/X _08789_/Y VGND VGND VPWR VPWR _09884_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11910_ _11909_/Y _11844_/X _11867_/Y VGND VGND VPWR VPWR _11910_/X sky130_fd_sc_hd__o21a_1
X_12890_ _12847_/X _12889_/Y _12847_/X _12889_/Y VGND VGND VPWR VPWR _12934_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11841_/A _11841_/B VGND VGND VPWR VPWR _11841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _15264_/A VGND VGND VPWR VPWR _14576_/A sky130_fd_sc_hd__buf_1
X_11772_ _12767_/A _11772_/B VGND VGND VPWR VPWR _11772_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13513_/A VGND VGND VPWR VPWR _15040_/A sky130_fd_sc_hd__buf_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10723_ _10723_/A VGND VGND VPWR VPWR _10723_/Y sky130_fd_sc_hd__inv_2
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14491_ _14464_/X _14490_/Y _14464_/X _14490_/Y VGND VGND VPWR VPWR _14516_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16230_ _16251_/B VGND VGND VPWR VPWR _16231_/B sky130_fd_sc_hd__buf_1
X_13442_ _13442_/A _13442_/B VGND VGND VPWR VPWR _13442_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10654_ _10654_/A _10654_/B VGND VGND VPWR VPWR _10654_/Y sky130_fd_sc_hd__nor2_1
X_16161_ _16268_/B VGND VGND VPWR VPWR _16334_/A sky130_fd_sc_hd__buf_1
X_13373_ _13313_/A _13313_/B _13313_/X _13372_/X VGND VGND VPWR VPWR _13373_/X sky130_fd_sc_hd__o22a_1
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10585_ _09970_/Y _10584_/A _09970_/A _10584_/Y _10940_/A VGND VGND VPWR VPWR _11904_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_127_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12324_ _12237_/X _12323_/Y _12237_/X _12323_/Y VGND VGND VPWR VPWR _12600_/A sky130_fd_sc_hd__a2bb2o_1
X_15112_ _15098_/X _15111_/Y _15098_/X _15111_/Y VGND VGND VPWR VPWR _15113_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16092_ _16032_/A _16032_/B _16032_/Y VGND VGND VPWR VPWR _16092_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12255_ _12255_/A VGND VGND VPWR VPWR _12255_/Y sky130_fd_sc_hd__inv_2
X_15043_ _15061_/A _15041_/X _15042_/X VGND VGND VPWR VPWR _15043_/X sky130_fd_sc_hd__o21a_1
X_11206_ _14056_/A _11206_/B VGND VGND VPWR VPWR _11206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12186_ _12166_/X _12185_/X _12166_/X _12185_/X VGND VGND VPWR VPWR _12257_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11137_ _12172_/A VGND VGND VPWR VPWR _12087_/A sky130_fd_sc_hd__inv_2
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15945_ _15948_/A _15948_/B VGND VGND VPWR VPWR _16023_/A sky130_fd_sc_hd__and2_1
XFILLER_95_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11068_ _12914_/A VGND VGND VPWR VPWR _12135_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15876_ _14220_/X _15842_/X _14220_/X _15842_/X VGND VGND VPWR VPWR _15890_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10019_ _08935_/A _09069_/A _08917_/A _08935_/X VGND VGND VPWR VPWR _10019_/X sky130_fd_sc_hd__a22o_1
X_14827_ _14774_/A _14774_/B _14774_/X _14826_/X VGND VGND VPWR VPWR _14827_/X sky130_fd_sc_hd__o22a_1
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14758_ _14757_/A _14757_/B _14757_/Y VGND VGND VPWR VPWR _14758_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14689_ _14663_/X _14688_/Y _14663_/X _14688_/Y VGND VGND VPWR VPWR _14741_/B sky130_fd_sc_hd__a2bb2o_1
X_13709_ _13709_/A VGND VGND VPWR VPWR _13709_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16428_ _16470_/Q VGND VGND VPWR VPWR _16428_/Y sky130_fd_sc_hd__inv_2
X_16359_ _16330_/A _16330_/B _16330_/Y VGND VGND VPWR VPWR _16359_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09802_ _09802_/A _09844_/A VGND VGND VPWR VPWR _09803_/B sky130_fd_sc_hd__or2_1
X_09733_ _09733_/A _09733_/B VGND VGND VPWR VPWR _09736_/A sky130_fd_sc_hd__or2_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09664_ _09995_/A _09664_/B VGND VGND VPWR VPWR _09664_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08615_ _09457_/B VGND VGND VPWR VPWR _09547_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09595_ _09595_/A _09595_/B VGND VGND VPWR VPWR _09595_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08546_ _08546_/A VGND VGND VPWR VPWR _08546_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08477_ input29/X input13/X VGND VGND VPWR VPWR _08477_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10370_ _10369_/Y _10309_/Y _10307_/Y VGND VGND VPWR VPWR _10370_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09029_ _09029_/A _09540_/B VGND VGND VPWR VPWR _09030_/B sky130_fd_sc_hd__or2_1
X_12040_ _13829_/A _12049_/B VGND VGND VPWR VPWR _12040_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13991_ _14832_/A _13991_/B VGND VGND VPWR VPWR _13991_/Y sky130_fd_sc_hd__nor2_1
X_15730_ _15682_/X _15729_/Y _15682_/X _15729_/Y VGND VGND VPWR VPWR _15815_/B sky130_fd_sc_hd__a2bb2o_1
X_12942_ _12942_/A _12942_/B VGND VGND VPWR VPWR _12942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15661_ _15661_/A VGND VGND VPWR VPWR _15947_/A sky130_fd_sc_hd__inv_2
XFILLER_65_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14612_ _14588_/A _14588_/B _14588_/Y VGND VGND VPWR VPWR _14612_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12873_ _12856_/A _12856_/B _12856_/Y VGND VGND VPWR VPWR _12873_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15592_ _15683_/A _15683_/B VGND VGND VPWR VPWR _15592_/Y sky130_fd_sc_hd__nor2_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _13621_/A _11839_/B VGND VGND VPWR VPWR _11824_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14543_ _14586_/A _14586_/B VGND VGND VPWR VPWR _14543_/Y sky130_fd_sc_hd__nor2_1
X_11755_ _11755_/A VGND VGND VPWR VPWR _11798_/A sky130_fd_sc_hd__inv_2
XFILLER_14_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14474_ _14474_/A _14474_/B VGND VGND VPWR VPWR _14474_/Y sky130_fd_sc_hd__nor2_1
X_10706_ _09653_/X _10705_/X _09653_/X _10705_/X VGND VGND VPWR VPWR _10707_/B sky130_fd_sc_hd__a2bb2oi_1
X_16213_ _16213_/A VGND VGND VPWR VPWR _16213_/Y sky130_fd_sc_hd__inv_2
X_13425_ _13359_/X _13424_/X _13359_/X _13424_/X VGND VGND VPWR VPWR _13425_/Y sky130_fd_sc_hd__a2bb2oi_1
X_11686_ _11657_/X _11685_/Y _11659_/B VGND VGND VPWR VPWR _11686_/X sky130_fd_sc_hd__o21a_1
X_10637_ _10637_/A VGND VGND VPWR VPWR _10637_/Y sky130_fd_sc_hd__inv_2
X_16144_ _16160_/A _16144_/B VGND VGND VPWR VPWR _16272_/A sky130_fd_sc_hd__or2_1
XFILLER_115_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13356_ _13350_/Y _13403_/A _13355_/X VGND VGND VPWR VPWR _13356_/Y sky130_fd_sc_hd__o21ai_1
X_10568_ _09275_/B _10244_/B _10244_/X VGND VGND VPWR VPWR _10569_/B sky130_fd_sc_hd__a21boi_1
X_16075_ _16039_/X _16074_/Y _16039_/X _16074_/Y VGND VGND VPWR VPWR _16108_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12307_ _14018_/A _12209_/B _12209_/Y VGND VGND VPWR VPWR _12307_/Y sky130_fd_sc_hd__o21ai_1
X_13287_ _13287_/A VGND VGND VPWR VPWR _13287_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10499_ _10499_/A VGND VGND VPWR VPWR _10499_/Y sky130_fd_sc_hd__inv_2
X_12238_ _13349_/A _12230_/B _12230_/Y _12237_/X VGND VGND VPWR VPWR _12238_/X sky130_fd_sc_hd__a2bb2o_1
X_15026_ _15028_/A _15028_/B VGND VGND VPWR VPWR _15082_/A sky130_fd_sc_hd__and2_1
XFILLER_123_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12169_ _12167_/A _12167_/B _12167_/X _12168_/Y VGND VGND VPWR VPWR _12261_/B sky130_fd_sc_hd__a22o_1
XFILLER_96_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15928_ _15896_/A _15896_/B _15896_/Y VGND VGND VPWR VPWR _15928_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 wbs_adr_i[12] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_2
XFILLER_76_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15859_ _15902_/A _15902_/B VGND VGND VPWR VPWR _15859_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08400_ _08662_/B _08400_/B VGND VGND VPWR VPWR _09677_/B sky130_fd_sc_hd__or2_1
XFILLER_64_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09380_ _09380_/A VGND VGND VPWR VPWR _09432_/B sky130_fd_sc_hd__inv_2
X_08331_ _08331_/A input32/X VGND VGND VPWR VPWR _08332_/B sky130_fd_sc_hd__nor2_1
X_08262_ input30/X VGND VGND VPWR VPWR _08263_/A sky130_fd_sc_hd__inv_2
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09716_ _09716_/A _09717_/B VGND VGND VPWR VPWR _10595_/A sky130_fd_sc_hd__and2_1
XFILLER_83_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09647_ _09975_/A _09650_/B VGND VGND VPWR VPWR _09647_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09558_/X _09577_/X _09558_/X _09577_/X VGND VGND VPWR VPWR _09664_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08529_ _08701_/A _08529_/B VGND VGND VPWR VPWR _09527_/A sky130_fd_sc_hd__or2_2
XFILLER_129_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11540_ _12440_/A _11631_/B VGND VGND VPWR VPWR _11540_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11471_ _12404_/A VGND VGND VPWR VPWR _14066_/A sky130_fd_sc_hd__buf_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14190_ _14190_/A _12631_/X VGND VGND VPWR VPWR _14190_/X sky130_fd_sc_hd__or2b_1
X_13210_ _14934_/A _13452_/B _13209_/Y VGND VGND VPWR VPWR _13210_/Y sky130_fd_sc_hd__o21ai_1
X_10422_ _10422_/A VGND VGND VPWR VPWR _10426_/A sky130_fd_sc_hd__inv_2
XFILLER_109_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13141_ _15234_/A VGND VGND VPWR VPWR _14953_/A sky130_fd_sc_hd__buf_1
X_10353_ _10423_/A VGND VGND VPWR VPWR _10421_/B sky130_fd_sc_hd__buf_1
X_13072_ _15252_/A _13113_/B VGND VGND VPWR VPWR _13072_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12023_ _12057_/A VGND VGND VPWR VPWR _13192_/A sky130_fd_sc_hd__buf_1
X_10284_ _13479_/B VGND VGND VPWR VPWR _10284_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15713_ _15550_/A _14926_/B _14926_/Y VGND VGND VPWR VPWR _15713_/X sky130_fd_sc_hd__o21a_1
X_13974_ _13973_/A _13973_/B _13973_/Y VGND VGND VPWR VPWR _13974_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12925_ _12911_/Y _12922_/Y _12924_/Y VGND VGND VPWR VPWR _12925_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15644_ _15644_/A _14380_/X VGND VGND VPWR VPWR _15644_/X sky130_fd_sc_hd__or2b_1
XFILLER_73_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12856_ _12856_/A _12856_/B VGND VGND VPWR VPWR _12856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15575_ _15700_/A _15575_/B VGND VGND VPWR VPWR _16055_/A sky130_fd_sc_hd__or2_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11807_/A VGND VGND VPWR VPWR _11854_/B sky130_fd_sc_hd__inv_2
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14474_/A _14474_/B _14471_/X _14474_/Y VGND VGND VPWR VPWR _14526_/X sky130_fd_sc_hd__o2bb2a_1
X_12787_ _12723_/Y _12786_/X _12723_/Y _12786_/X VGND VGND VPWR VPWR _12788_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11738_ _11742_/B _11737_/Y _11742_/B _11737_/Y VGND VGND VPWR VPWR _11777_/B sky130_fd_sc_hd__o2bb2a_1
X_11669_ _11668_/A _15433_/A _11668_/Y VGND VGND VPWR VPWR _11669_/X sky130_fd_sc_hd__a21o_1
X_14457_ _14459_/A _14459_/B VGND VGND VPWR VPWR _14457_/Y sky130_fd_sc_hd__nor2_1
X_14388_ _14388_/A _15958_/A VGND VGND VPWR VPWR _14388_/X sky130_fd_sc_hd__or2_1
X_13408_ _14901_/A _13408_/B VGND VGND VPWR VPWR _13408_/X sky130_fd_sc_hd__and2_1
XFILLER_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16127_ _15992_/A _16056_/X _15991_/X VGND VGND VPWR VPWR _16127_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13339_ _13278_/A _13338_/Y _13278_/A _13338_/Y VGND VGND VPWR VPWR _13340_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16058_ _16125_/A _16125_/B VGND VGND VPWR VPWR _16058_/X sky130_fd_sc_hd__and2_1
X_15009_ _12088_/X _15005_/X _12088_/X _15005_/X VGND VGND VPWR VPWR _15044_/B sky130_fd_sc_hd__a2bb2o_1
X_08880_ _08982_/A _08982_/B VGND VGND VPWR VPWR _08880_/X sky130_fd_sc_hd__and2_1
XFILLER_69_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09501_ _08839_/A _09461_/X _08839_/A _09461_/X VGND VGND VPWR VPWR _09502_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09432_ _09432_/A _09432_/B VGND VGND VPWR VPWR _09432_/X sky130_fd_sc_hd__or2_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09363_ _09363_/A VGND VGND VPWR VPWR _09429_/B sky130_fd_sc_hd__inv_2
XFILLER_40_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08314_ _08314_/A VGND VGND VPWR VPWR _08314_/Y sky130_fd_sc_hd__inv_2
X_09294_ _09293_/A _09293_/B _08929_/A _09293_/Y VGND VGND VPWR VPWR _09298_/B sky130_fd_sc_hd__o2bb2a_1
X_08245_ input5/X _08245_/B VGND VGND VPWR VPWR _08312_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10971_ _10241_/B _10151_/B _10151_/Y VGND VGND VPWR VPWR _10972_/A sky130_fd_sc_hd__a21oi_1
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13690_ _13676_/Y _13688_/X _13689_/Y VGND VGND VPWR VPWR _13690_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12710_ _12703_/A _12703_/B _12703_/X _12709_/X VGND VGND VPWR VPWR _12710_/X sky130_fd_sc_hd__o22a_1
X_12641_ _12641_/A VGND VGND VPWR VPWR _12641_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12572_ _12569_/Y _12571_/Y _12569_/A _12571_/A _12501_/A VGND VGND VPWR VPWR _12623_/B
+ sky130_fd_sc_hd__o221a_1
X_15360_ _15360_/A _15351_/X VGND VGND VPWR VPWR _15360_/X sky130_fd_sc_hd__or2b_1
XFILLER_11_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14311_ _14274_/A _14310_/Y _14274_/A _14310_/Y VGND VGND VPWR VPWR _14394_/B sky130_fd_sc_hd__a2bb2o_1
X_15291_ _15234_/A _15234_/B _15234_/Y VGND VGND VPWR VPWR _15291_/Y sky130_fd_sc_hd__o21ai_1
X_11523_ _11528_/A VGND VGND VPWR VPWR _11612_/A sky130_fd_sc_hd__inv_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14242_ _14243_/A _14243_/B VGND VGND VPWR VPWR _14372_/A sky130_fd_sc_hd__and2_1
X_11454_ _11448_/Y _12544_/A _11453_/Y VGND VGND VPWR VPWR _12538_/A sky130_fd_sc_hd__o21ai_1
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10405_ _10405_/A VGND VGND VPWR VPWR _11780_/A sky130_fd_sc_hd__buf_1
XFILLER_124_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14173_ _15910_/A _14288_/B VGND VGND VPWR VPWR _14295_/A sky130_fd_sc_hd__and2_1
X_11385_ _08907_/X _11385_/B VGND VGND VPWR VPWR _11385_/X sky130_fd_sc_hd__and2b_1
XFILLER_112_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13124_ _13047_/Y _13122_/X _13123_/Y VGND VGND VPWR VPWR _13124_/X sky130_fd_sc_hd__o21a_1
X_10336_ _11724_/A _10335_/B _10335_/Y VGND VGND VPWR VPWR _10336_/Y sky130_fd_sc_hd__a21oi_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13055_ _13055_/A _13028_/X VGND VGND VPWR VPWR _13055_/X sky130_fd_sc_hd__or2b_1
X_10267_ _10288_/B VGND VGND VPWR VPWR _10268_/A sky130_fd_sc_hd__inv_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ _13641_/A _12071_/B _12005_/Y VGND VGND VPWR VPWR _12006_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10198_ _10197_/Y _10134_/X _10197_/Y _10134_/X VGND VGND VPWR VPWR _10198_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13957_ _13901_/Y _13955_/X _13956_/Y VGND VGND VPWR VPWR _13957_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12908_ _13609_/A VGND VGND VPWR VPWR _12923_/A sky130_fd_sc_hd__buf_1
XFILLER_62_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15627_ _16036_/A VGND VGND VPWR VPWR _15673_/A sky130_fd_sc_hd__inv_2
X_13888_ _13861_/X _13887_/Y _13861_/X _13887_/Y VGND VGND VPWR VPWR _13962_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12839_ _12825_/Y _12837_/X _12838_/Y VGND VGND VPWR VPWR _12839_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _15555_/X _15557_/Y _15555_/X _15557_/Y VGND VGND VPWR VPWR _15558_/X sky130_fd_sc_hd__a2bb2o_1
X_15489_ _15437_/A _15437_/B _15437_/A _15437_/B VGND VGND VPWR VPWR _15489_/X sky130_fd_sc_hd__a2bb2o_1
X_14509_ _15216_/A _14508_/B _13007_/Y _14508_/Y VGND VGND VPWR VPWR _14509_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 wbs_dat_i[6] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__buf_1
XFILLER_115_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09981_ _09981_/A _09981_/B VGND VGND VPWR VPWR _09981_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08932_ _10228_/B _08932_/B VGND VGND VPWR VPWR _08932_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08863_ _08795_/X _08801_/A _08803_/Y _08862_/X VGND VGND VPWR VPWR _08863_/X sky130_fd_sc_hd__o22a_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08794_ _08794_/A VGND VGND VPWR VPWR _09492_/A sky130_fd_sc_hd__buf_1
XFILLER_29_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09415_ _09415_/A _09415_/B VGND VGND VPWR VPWR _09415_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09346_ _09561_/A _09346_/B VGND VGND VPWR VPWR _09347_/A sky130_fd_sc_hd__or2_1
X_09277_ _09241_/X _09276_/X _09241_/X _09276_/X VGND VGND VPWR VPWR _10438_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_32_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11170_ _13048_/A _11170_/B VGND VGND VPWR VPWR _11170_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10121_ _10120_/X _08989_/Y _10120_/X _08989_/Y VGND VGND VPWR VPWR _10237_/B sky130_fd_sc_hd__a2bb2o_1
X_10052_ _10052_/A _10077_/B VGND VGND VPWR VPWR _10052_/X sky130_fd_sc_hd__and2_1
XFILLER_102_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14860_ _14829_/X _14859_/X _14829_/X _14859_/X VGND VGND VPWR VPWR _14930_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14791_ _15455_/A VGND VGND VPWR VPWR _14794_/A sky130_fd_sc_hd__buf_1
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13811_ _13768_/X _13810_/X _13768_/X _13810_/X VGND VGND VPWR VPWR _13852_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13742_ _14493_/A _13691_/B _13691_/Y VGND VGND VPWR VPWR _13742_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_90_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10954_ _13510_/A _10953_/B _10953_/X _10802_/X VGND VGND VPWR VPWR _10954_/X sky130_fd_sc_hd__o22a_1
XFILLER_43_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16461_ _16357_/A _16461_/D VGND VGND VPWR VPWR _16461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13673_ _14493_/A _13691_/B VGND VGND VPWR VPWR _13673_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10885_ _10885_/A VGND VGND VPWR VPWR _10885_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16392_ _16392_/A _16392_/B _16392_/C VGND VGND VPWR VPWR _16454_/A sky130_fd_sc_hd__or3_1
X_12624_ _14214_/A _12622_/X _12623_/X VGND VGND VPWR VPWR _12624_/X sky130_fd_sc_hd__o21a_1
X_15412_ _15412_/A _15412_/B VGND VGND VPWR VPWR _15412_/X sky130_fd_sc_hd__or2_1
X_12555_ _15534_/A VGND VGND VPWR VPWR _14914_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15343_ _15343_/A _15343_/B VGND VGND VPWR VPWR _15343_/X sky130_fd_sc_hd__or2_1
XFILLER_8_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11506_ _11506_/A VGND VGND VPWR VPWR _13501_/A sky130_fd_sc_hd__buf_1
XFILLER_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12486_ _12486_/A _12486_/B VGND VGND VPWR VPWR _12486_/Y sky130_fd_sc_hd__nand2_1
X_15274_ _14576_/A _15264_/B _15264_/Y _15273_/Y VGND VGND VPWR VPWR _15274_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14225_ _14231_/A _14225_/B VGND VGND VPWR VPWR _15878_/A sky130_fd_sc_hd__or2_1
X_11437_ _14032_/A _11224_/B _11224_/Y VGND VGND VPWR VPWR _11437_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11368_ _14060_/A _11188_/B _11188_/Y VGND VGND VPWR VPWR _11368_/Y sky130_fd_sc_hd__o21ai_1
X_14156_ _14075_/X _14155_/Y _14075_/X _14155_/Y VGND VGND VPWR VPWR _14245_/A sky130_fd_sc_hd__a2bb2o_4
X_13107_ _15261_/A _13107_/B VGND VGND VPWR VPWR _13107_/Y sky130_fd_sc_hd__nand2_1
X_10319_ _13525_/A _10319_/B VGND VGND VPWR VPWR _10319_/X sky130_fd_sc_hd__and2_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14087_ _14901_/A _14084_/B _14084_/X _14086_/Y VGND VGND VPWR VPWR _14091_/B sky130_fd_sc_hd__o22a_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11299_ _11297_/Y _11298_/Y _11298_/B _09926_/X _10792_/X VGND VGND VPWR VPWR _12944_/A
+ sky130_fd_sc_hd__o221a_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13883_/A VGND VGND VPWR VPWR _15234_/A sky130_fd_sc_hd__buf_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14989_ _14956_/A _14956_/B _14956_/Y _14959_/X VGND VGND VPWR VPWR _14989_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09200_ _09196_/Y _09199_/A _09198_/X _09199_/Y VGND VGND VPWR VPWR _09200_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09131_ _09424_/A _09131_/B VGND VGND VPWR VPWR _09131_/Y sky130_fd_sc_hd__nand2_1
X_09062_ _08831_/X _09043_/Y _08831_/X _09043_/Y VGND VGND VPWR VPWR _10018_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09964_ _09997_/A _09997_/B VGND VGND VPWR VPWR _09964_/X sky130_fd_sc_hd__and2_1
XFILLER_131_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _09883_/A _09883_/B _09884_/B VGND VGND VPWR VPWR _09903_/A sky130_fd_sc_hd__a21bo_1
X_08915_ _09401_/A VGND VGND VPWR VPWR _09817_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _09826_/B VGND VGND VPWR VPWR _08847_/A sky130_fd_sc_hd__inv_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08777_ _10011_/A VGND VGND VPWR VPWR _08778_/A sky130_fd_sc_hd__buf_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10670_ _11918_/A VGND VGND VPWR VPWR _11859_/A sky130_fd_sc_hd__inv_2
XFILLER_41_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09329_ _09328_/A _09328_/B _09328_/X VGND VGND VPWR VPWR _09330_/B sky130_fd_sc_hd__a21boi_1
XFILLER_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12340_ _12336_/Y _12569_/A _12339_/Y VGND VGND VPWR VPWR _12344_/B sky130_fd_sc_hd__o21ai_2
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12271_ _11326_/A _12270_/A _11326_/Y _12270_/Y VGND VGND VPWR VPWR _12273_/B sky130_fd_sc_hd__o22a_1
XFILLER_107_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14010_ _15416_/A _13958_/B _13958_/Y VGND VGND VPWR VPWR _14010_/Y sky130_fd_sc_hd__o21ai_1
X_11222_ _11222_/A _11083_/X VGND VGND VPWR VPWR _11222_/X sky130_fd_sc_hd__or2b_1
XFILLER_4_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11153_ _11141_/X _11152_/Y _11141_/X _11152_/Y VGND VGND VPWR VPWR _11312_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15961_ _16005_/A _15959_/X _15960_/X VGND VGND VPWR VPWR _15961_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11084_ _11222_/A _11082_/X _11083_/X VGND VGND VPWR VPWR _11084_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10104_ _10103_/A _10103_/B _10123_/B VGND VGND VPWR VPWR _10177_/A sky130_fd_sc_hd__o21ai_2
X_14912_ _14912_/A _14912_/B VGND VGND VPWR VPWR _14912_/Y sky130_fd_sc_hd__nand2_1
X_15892_ _15892_/A _15892_/B VGND VGND VPWR VPWR _15892_/Y sky130_fd_sc_hd__nand2_1
X_10035_ _10035_/A _10035_/B VGND VGND VPWR VPWR _10035_/Y sky130_fd_sc_hd__nor2_1
X_14843_ _14838_/X _14842_/X _14838_/X _14842_/X VGND VGND VPWR VPWR _14944_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14774_ _14774_/A _14774_/B VGND VGND VPWR VPWR _14774_/X sky130_fd_sc_hd__and2_1
XFILLER_90_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11986_ _11986_/A VGND VGND VPWR VPWR _11986_/Y sky130_fd_sc_hd__inv_2
X_13725_ _13702_/X _13724_/X _13702_/X _13724_/X VGND VGND VPWR VPWR _13773_/B sky130_fd_sc_hd__a2bb2o_1
X_10937_ _10935_/Y _10936_/Y _10839_/Y VGND VGND VPWR VPWR _11116_/A sky130_fd_sc_hd__o21ai_2
X_16444_ _16434_/A _16434_/B _16434_/Y _16439_/X _16443_/Y VGND VGND VPWR VPWR _16444_/Y
+ sky130_fd_sc_hd__a2111oi_2
X_13656_ _15122_/A _13642_/B _13642_/Y VGND VGND VPWR VPWR _13656_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12607_ _14244_/A _12607_/B VGND VGND VPWR VPWR _12607_/Y sky130_fd_sc_hd__nand2_1
X_10868_ _09415_/A _09415_/B _09415_/Y VGND VGND VPWR VPWR _10869_/A sky130_fd_sc_hd__o21ai_1
X_16375_ _16320_/A _16320_/B _16320_/Y VGND VGND VPWR VPWR _16375_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13587_ _13641_/A _13642_/B VGND VGND VPWR VPWR _13587_/Y sky130_fd_sc_hd__nor2_1
X_10799_ _10798_/A _10798_/B _10798_/Y _09393_/A VGND VGND VPWR VPWR _10951_/A sky130_fd_sc_hd__o211a_1
X_12538_ _12538_/A _12538_/B VGND VGND VPWR VPWR _12538_/Y sky130_fd_sc_hd__nand2_1
X_15326_ _15331_/A _15331_/B VGND VGND VPWR VPWR _15326_/Y sky130_fd_sc_hd__nor2_1
X_15257_ _15220_/X _15256_/Y _15220_/X _15256_/Y VGND VGND VPWR VPWR _15258_/B sky130_fd_sc_hd__a2bb2o_1
X_12469_ _12461_/Y _12468_/X _12461_/Y _12468_/X VGND VGND VPWR VPWR _12469_/Y sky130_fd_sc_hd__a2bb2oi_1
X_14208_ _14208_/A _12625_/X VGND VGND VPWR VPWR _14208_/X sky130_fd_sc_hd__or2b_1
XFILLER_125_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15188_ _15122_/A _15122_/B _15122_/Y VGND VGND VPWR VPWR _15188_/Y sky130_fd_sc_hd__o21ai_1
X_14139_ _14139_/A VGND VGND VPWR VPWR _14139_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ _08239_/Y _08699_/A _08239_/A _08699_/Y VGND VGND VPWR VPWR _08701_/B sky130_fd_sc_hd__o22a_1
X_09680_ _09680_/A _09829_/B VGND VGND VPWR VPWR _09683_/A sky130_fd_sc_hd__or2_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08631_ _09225_/B VGND VGND VPWR VPWR _08631_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08562_ _08561_/A _08333_/Y _08561_/Y _08333_/A VGND VGND VPWR VPWR _08563_/B sky130_fd_sc_hd__o22a_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08493_ _08316_/A _08248_/B _08471_/Y _08527_/A VGND VGND VPWR VPWR _08516_/A sky130_fd_sc_hd__o22a_1
XFILLER_62_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09114_ _09110_/Y _09112_/Y _09113_/Y VGND VGND VPWR VPWR _09118_/B sky130_fd_sc_hd__o21ai_1
X_09045_ _08716_/A _08716_/B _08716_/X _09044_/X VGND VGND VPWR VPWR _09045_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09947_ _09947_/A VGND VGND VPWR VPWR _09947_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09868_/X _08781_/Y _09868_/X _08781_/Y VGND VGND VPWR VPWR _09885_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08829_ _09225_/A _09457_/B _08717_/X VGND VGND VPWR VPWR _08830_/A sky130_fd_sc_hd__o21ai_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11840_ _11824_/Y _11838_/X _11839_/Y VGND VGND VPWR VPWR _11840_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11771_/A VGND VGND VPWR VPWR _12767_/A sky130_fd_sc_hd__buf_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13510_ _13510_/A _13510_/B VGND VGND VPWR VPWR _13510_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10722_ _10722_/A VGND VGND VPWR VPWR _10722_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14490_ _14465_/A _14465_/B _14465_/Y VGND VGND VPWR VPWR _14490_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13441_ _13390_/Y _13439_/X _13440_/Y VGND VGND VPWR VPWR _13441_/X sky130_fd_sc_hd__o21a_1
X_10653_ _10653_/A VGND VGND VPWR VPWR _10653_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16160_ _16160_/A _16160_/B VGND VGND VPWR VPWR _16268_/B sky130_fd_sc_hd__or2_1
X_13372_ _13379_/A _13370_/X _13371_/X VGND VGND VPWR VPWR _13372_/X sky130_fd_sc_hd__o21a_1
X_10584_ _10584_/A VGND VGND VPWR VPWR _10584_/Y sky130_fd_sc_hd__inv_2
X_16091_ _16094_/A _16094_/B VGND VGND VPWR VPWR _16091_/Y sky130_fd_sc_hd__nor2_1
X_12323_ _12230_/A _12230_/B _12230_/Y VGND VGND VPWR VPWR _12323_/Y sky130_fd_sc_hd__o21ai_1
X_15111_ _15054_/A _15054_/B _15054_/Y VGND VGND VPWR VPWR _15111_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15042_ _15042_/A _15042_/B VGND VGND VPWR VPWR _15042_/X sky130_fd_sc_hd__or2_1
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12254_ _12254_/A _12254_/B VGND VGND VPWR VPWR _12254_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11205_ _11088_/X _11204_/X _11088_/X _11204_/X VGND VGND VPWR VPWR _11206_/B sky130_fd_sc_hd__a2bb2o_1
X_12185_ _13713_/A _12259_/B _12259_/A _12259_/B VGND VGND VPWR VPWR _12185_/X sky130_fd_sc_hd__a2bb2o_1
X_11136_ _11138_/A VGND VGND VPWR VPWR _11136_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15944_ _15885_/X _15943_/Y _15885_/X _15943_/Y VGND VGND VPWR VPWR _15948_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11067_ _12826_/A VGND VGND VPWR VPWR _12914_/A sky130_fd_sc_hd__buf_1
XFILLER_49_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15875_ _15875_/A VGND VGND VPWR VPWR _15890_/A sky130_fd_sc_hd__inv_2
XFILLER_49_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10018_ _10018_/A _10018_/B VGND VGND VPWR VPWR _10061_/B sky130_fd_sc_hd__nor2_1
X_14826_ _14778_/A _14778_/B _14778_/X _14825_/X VGND VGND VPWR VPWR _14826_/X sky130_fd_sc_hd__o22a_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14757_ _14757_/A _14757_/B VGND VGND VPWR VPWR _14757_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11969_ _11951_/Y _11967_/X _11968_/Y VGND VGND VPWR VPWR _11969_/X sky130_fd_sc_hd__o21a_1
X_13708_ _13716_/A VGND VGND VPWR VPWR _15116_/A sky130_fd_sc_hd__buf_1
X_14688_ _15349_/A _14743_/B _14687_/Y VGND VGND VPWR VPWR _14688_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16427_ _16412_/Y _16415_/X _16416_/Y _16420_/X _16426_/X VGND VGND VPWR VPWR _16445_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13639_ _13590_/Y _13636_/Y _13638_/Y VGND VGND VPWR VPWR _13640_/A sky130_fd_sc_hd__o21ai_1
XFILLER_20_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16358_ _16358_/A VGND VGND VPWR VPWR _16358_/X sky130_fd_sc_hd__buf_1
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15309_ _14584_/A _15252_/B _15252_/Y VGND VGND VPWR VPWR _15309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16289_ _16265_/X _16288_/Y _16265_/X _16288_/Y VGND VGND VPWR VPWR _16332_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09801_ _09801_/A _09801_/B VGND VGND VPWR VPWR _09844_/A sky130_fd_sc_hd__or2_1
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09732_ _08567_/X _09734_/B _08567_/X _09734_/B VGND VGND VPWR VPWR _09733_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09663_ _09585_/Y _09661_/X _09662_/Y VGND VGND VPWR VPWR _09663_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08614_ _08650_/A _08614_/B VGND VGND VPWR VPWR _09457_/B sky130_fd_sc_hd__or2_1
X_09594_ _09986_/A VGND VGND VPWR VPWR _09987_/A sky130_fd_sc_hd__buf_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _09740_/A _08567_/B VGND VGND VPWR VPWR _08546_/A sky130_fd_sc_hd__or2_1
X_08476_ input30/X input14/X VGND VGND VPWR VPWR _08476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09028_ _09028_/A VGND VGND VPWR VPWR _09540_/B sky130_fd_sc_hd__inv_2
XFILLER_2_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13990_ _14956_/A _13989_/B _13989_/Y VGND VGND VPWR VPWR _13990_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12941_ _12879_/Y _12939_/X _12940_/Y VGND VGND VPWR VPWR _12941_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15660_ _16027_/A VGND VGND VPWR VPWR _15665_/A sky130_fd_sc_hd__inv_2
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12872_ _12942_/A VGND VGND VPWR VPWR _14677_/A sky130_fd_sc_hd__buf_1
XFILLER_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14611_ _14611_/A VGND VGND VPWR VPWR _15345_/A sky130_fd_sc_hd__buf_1
XFILLER_73_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11823_ _11795_/X _11822_/X _11795_/X _11822_/X VGND VGND VPWR VPWR _11839_/B sky130_fd_sc_hd__a2bb2o_1
X_15591_ _14393_/X _15590_/X _14393_/X _15590_/X VGND VGND VPWR VPWR _15683_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14521_/X _14541_/X _14521_/X _14541_/X VGND VGND VPWR VPWR _14586_/B sky130_fd_sc_hd__a2bb2o_1
X_11754_ _11771_/A _11741_/B _11741_/X _11753_/Y VGND VGND VPWR VPWR _11798_/B sky130_fd_sc_hd__a22o_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11685_/A VGND VGND VPWR VPWR _11685_/Y sky130_fd_sc_hd__inv_2
X_14473_ _11929_/Y _14472_/X _11929_/Y _14472_/X VGND VGND VPWR VPWR _14474_/B sky130_fd_sc_hd__o2bb2a_1
X_10705_ _09981_/A _09654_/B _09654_/Y VGND VGND VPWR VPWR _10705_/X sky130_fd_sc_hd__o21a_1
X_16212_ _16094_/A _16094_/B _16094_/Y VGND VGND VPWR VPWR _16214_/A sky130_fd_sc_hd__o21ai_1
X_13424_ _13337_/A _13337_/B _13337_/A _13337_/B VGND VGND VPWR VPWR _13424_/X sky130_fd_sc_hd__a2bb2o_1
X_10636_ _10600_/Y _10634_/Y _10635_/Y VGND VGND VPWR VPWR _10637_/A sky130_fd_sc_hd__o21ai_1
X_16143_ _15820_/X _16142_/X _15820_/X _16142_/X VGND VGND VPWR VPWR _16144_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13355_ _15473_/A _13355_/B VGND VGND VPWR VPWR _13355_/X sky130_fd_sc_hd__or2_1
X_10567_ _10555_/X _10566_/Y _10555_/X _10566_/Y VGND VGND VPWR VPWR _10671_/A sky130_fd_sc_hd__o2bb2a_1
X_16074_ _16040_/A _16040_/B _16040_/Y VGND VGND VPWR VPWR _16074_/Y sky130_fd_sc_hd__o21ai_1
X_12306_ _12306_/A _12306_/B VGND VGND VPWR VPWR _12306_/Y sky130_fd_sc_hd__nand2_1
X_13286_ _13250_/Y _13284_/Y _13285_/Y VGND VGND VPWR VPWR _13287_/A sky130_fd_sc_hd__o21ai_1
X_10498_ _09838_/A _09838_/B _09839_/A VGND VGND VPWR VPWR _10499_/A sky130_fd_sc_hd__o21ai_1
X_12237_ _13351_/A _12236_/B _12235_/X _12236_/Y VGND VGND VPWR VPWR _12237_/X sky130_fd_sc_hd__a2bb2o_1
X_15025_ _11725_/Y _14997_/X _11725_/Y _14997_/X VGND VGND VPWR VPWR _15028_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12168_ _12168_/A VGND VGND VPWR VPWR _12168_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12099_ _13703_/A _12160_/B _12098_/Y VGND VGND VPWR VPWR _12099_/Y sky130_fd_sc_hd__o21ai_1
X_11119_ _11119_/A VGND VGND VPWR VPWR _11119_/Y sky130_fd_sc_hd__inv_2
X_15927_ _15960_/A _15960_/B VGND VGND VPWR VPWR _16005_/A sky130_fd_sc_hd__and2_1
XFILLER_110_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 wbs_adr_i[13] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15858_ _14184_/X _15848_/X _14184_/X _15848_/X VGND VGND VPWR VPWR _15902_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15789_ _15784_/Y _15786_/Y _15788_/Y VGND VGND VPWR VPWR _15794_/B sky130_fd_sc_hd__o21ai_1
X_14809_ _14809_/A _14809_/B VGND VGND VPWR VPWR _14809_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08330_ _08328_/Y _08329_/A _08328_/A _08329_/Y _08304_/A VGND VGND VPWR VPWR _08565_/B
+ sky130_fd_sc_hd__o221a_1
X_08261_ input14/X VGND VGND VPWR VPWR _08341_/B sky130_fd_sc_hd__inv_2
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09715_ _09409_/A _09713_/A _10216_/A _09714_/Y VGND VGND VPWR VPWR _09717_/B sky130_fd_sc_hd__o22a_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09646_ _09642_/Y _10731_/A _09645_/Y VGND VGND VPWR VPWR _09650_/B sky130_fd_sc_hd__o21ai_1
XFILLER_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _08692_/A _09154_/A _09528_/A VGND VGND VPWR VPWR _09577_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08527_/A _08318_/Y _08527_/Y _08318_/A VGND VGND VPWR VPWR _08529_/B sky130_fd_sc_hd__o22a_1
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08459_ _08459_/A VGND VGND VPWR VPWR _08459_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11470_ _13313_/A VGND VGND VPWR VPWR _12404_/A sky130_fd_sc_hd__inv_2
X_10421_ _10421_/A _10421_/B VGND VGND VPWR VPWR _10422_/A sky130_fd_sc_hd__or2_1
XFILLER_124_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13140_ _15289_/A _13139_/B _13139_/Y VGND VGND VPWR VPWR _13140_/X sky130_fd_sc_hd__a21o_1
X_10352_ _10352_/A _10620_/A VGND VGND VPWR VPWR _10423_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13071_ _13021_/X _13070_/X _13021_/X _13070_/X VGND VGND VPWR VPWR _13113_/B sky130_fd_sc_hd__a2bb2o_1
X_12022_ _13194_/A _12059_/B VGND VGND VPWR VPWR _12022_/Y sky130_fd_sc_hd__nor2_1
X_10283_ _10282_/A _11721_/A _10282_/Y _10206_/A VGND VGND VPWR VPWR _13479_/B sky130_fd_sc_hd__o22a_1
XFILLER_105_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13973_ _13973_/A _13973_/B VGND VGND VPWR VPWR _13973_/Y sky130_fd_sc_hd__nor2_1
X_15712_ _16123_/A _15821_/B VGND VGND VPWR VPWR _15712_/X sky130_fd_sc_hd__and2_1
XFILLER_74_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12924_ _14459_/A _12924_/B VGND VGND VPWR VPWR _12924_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15643_ _16032_/A VGND VGND VPWR VPWR _15669_/A sky130_fd_sc_hd__inv_2
X_12855_ _12801_/Y _12853_/X _12854_/Y VGND VGND VPWR VPWR _12855_/X sky130_fd_sc_hd__o21a_1
X_15574_ _15551_/X _15573_/X _15551_/X _15573_/X VGND VGND VPWR VPWR _15575_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12786_ _12726_/Y _12784_/X _12785_/Y VGND VGND VPWR VPWR _12786_/X sky130_fd_sc_hd__o21a_1
X_11806_ _10374_/A _11761_/A _10453_/B _11805_/Y VGND VGND VPWR VPWR _11807_/A sky130_fd_sc_hd__o22a_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14477_/A _14477_/B _14470_/X _14477_/Y VGND VGND VPWR VPWR _14525_/X sky130_fd_sc_hd__o2bb2a_1
X_11737_ _10325_/B _11743_/A _11736_/Y VGND VGND VPWR VPWR _11737_/Y sky130_fd_sc_hd__a21oi_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11668_ _11668_/A _12486_/A VGND VGND VPWR VPWR _11668_/Y sky130_fd_sc_hd__nor2_1
X_14456_ _14431_/X _14455_/X _14431_/X _14455_/X VGND VGND VPWR VPWR _14459_/B sky130_fd_sc_hd__a2bb2o_1
X_14387_ _15620_/A _14385_/X _14386_/X VGND VGND VPWR VPWR _14387_/X sky130_fd_sc_hd__o21a_1
X_13407_ _14904_/A _13405_/B _13405_/X _14240_/A VGND VGND VPWR VPWR _13408_/B sky130_fd_sc_hd__o22a_1
X_10619_ _15212_/A VGND VGND VPWR VPWR _11886_/A sky130_fd_sc_hd__inv_2
X_11599_ _11599_/A _11599_/B VGND VGND VPWR VPWR _11599_/Y sky130_fd_sc_hd__nand2_1
X_16126_ _16058_/X _16124_/X _16386_/B VGND VGND VPWR VPWR _16126_/Y sky130_fd_sc_hd__o21ai_1
X_13338_ _14727_/A _13279_/B _13279_/Y VGND VGND VPWR VPWR _13338_/Y sky130_fd_sc_hd__o21ai_1
X_16057_ _15992_/X _16056_/X _15992_/X _16056_/X VGND VGND VPWR VPWR _16125_/B sky130_fd_sc_hd__a2bb2o_1
X_13269_ _15087_/A VGND VGND VPWR VPWR _14722_/A sky130_fd_sc_hd__buf_1
X_15008_ _15046_/A _15046_/B VGND VGND VPWR VPWR _15055_/A sky130_fd_sc_hd__and2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09500_ _09500_/A _09500_/B VGND VGND VPWR VPWR _09500_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09431_ _09431_/A _09431_/B VGND VGND VPWR VPWR _09431_/X sky130_fd_sc_hd__or2_1
X_09362_ _09361_/X _09358_/X _09361_/X _09358_/X VGND VGND VPWR VPWR _09363_/A sky130_fd_sc_hd__a2bb2o_1
X_08313_ _08313_/A VGND VGND VPWR VPWR _08313_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09293_ _09293_/A _09293_/B VGND VGND VPWR VPWR _09293_/Y sky130_fd_sc_hd__nor2_1
X_08244_ input21/X VGND VGND VPWR VPWR _08245_/B sky130_fd_sc_hd__inv_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10970_ _10970_/A VGND VGND VPWR VPWR _12174_/A sky130_fd_sc_hd__inv_2
XFILLER_28_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09629_ _09629_/A _09629_/B _09707_/A VGND VGND VPWR VPWR _09629_/X sky130_fd_sc_hd__and3_1
X_12640_ _14171_/A _12638_/X _12639_/X VGND VGND VPWR VPWR _12641_/A sky130_fd_sc_hd__o21ai_1
XFILLER_70_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14310_ _15857_/A _14275_/B _14275_/Y VGND VGND VPWR VPWR _14310_/Y sky130_fd_sc_hd__o21ai_1
X_12571_ _12571_/A VGND VGND VPWR VPWR _12571_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15290_ _15289_/A _15289_/B _15289_/Y VGND VGND VPWR VPWR _15290_/X sky130_fd_sc_hd__a21o_1
X_11522_ _11604_/A _11522_/B VGND VGND VPWR VPWR _11528_/A sky130_fd_sc_hd__or2_1
X_14241_ _14240_/A _14239_/Y _14244_/B _14239_/A _14245_/A VGND VGND VPWR VPWR _14243_/B
+ sky130_fd_sc_hd__a221o_1
X_11453_ _15540_/A _11453_/B VGND VGND VPWR VPWR _11453_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14172_ _12638_/X _14171_/X _12638_/X _14171_/X VGND VGND VPWR VPWR _14288_/B sky130_fd_sc_hd__a2bb2o_1
X_10404_ _10402_/A _10403_/A _10402_/Y _10403_/Y _09392_/A VGND VGND VPWR VPWR _10405_/A
+ sky130_fd_sc_hd__o221a_1
X_11384_ _12312_/A _11384_/B VGND VGND VPWR VPWR _11384_/Y sky130_fd_sc_hd__nand2_1
X_13123_ _15237_/A _13123_/B VGND VGND VPWR VPWR _13123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10335_ _11724_/A _10335_/B VGND VGND VPWR VPWR _10335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13054_ _13773_/A VGND VGND VPWR VPWR _15243_/A sky130_fd_sc_hd__buf_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _09344_/X _10265_/X _09344_/X _10265_/X VGND VGND VPWR VPWR _10288_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12005_ _12005_/A _12071_/B VGND VGND VPWR VPWR _12005_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10197_ _10120_/X _08989_/Y _08468_/Y VGND VGND VPWR VPWR _10197_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_19_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13956_ _15414_/A _13956_/B VGND VGND VPWR VPWR _13956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13887_ _14832_/A _13991_/B _13886_/Y VGND VGND VPWR VPWR _13887_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12907_ _14461_/A _12926_/B VGND VGND VPWR VPWR _12907_/Y sky130_fd_sc_hd__nor2_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ _15624_/A _15625_/A _15624_/Y _15625_/Y _15571_/A VGND VGND VPWR VPWR _16036_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12838_ _15084_/A _12838_/B VGND VGND VPWR VPWR _12838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15556_/Y _15229_/Y _15174_/Y VGND VGND VPWR VPWR _15557_/Y sky130_fd_sc_hd__o21ai_1
X_12769_ _12769_/A _12769_/B VGND VGND VPWR VPWR _12769_/Y sky130_fd_sc_hd__nand2_1
X_15488_ _15554_/A _15554_/B VGND VGND VPWR VPWR _15488_/Y sky130_fd_sc_hd__nor2_1
X_14508_ _15216_/A _14508_/B VGND VGND VPWR VPWR _14508_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput20 wbs_dat_i[11] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_4
X_14439_ _14439_/A _14439_/B VGND VGND VPWR VPWR _14439_/Y sky130_fd_sc_hd__nor2_1
Xinput31 wbs_dat_i[7] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16109_ _16076_/X _16107_/X _16179_/B VGND VGND VPWR VPWR _16109_/X sky130_fd_sc_hd__o21a_1
X_09980_ _09980_/A _09981_/B VGND VGND VPWR VPWR _09980_/Y sky130_fd_sc_hd__nor2_1
X_08931_ _08931_/A VGND VGND VPWR VPWR _08931_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08862_ _09494_/A _08809_/Y _08810_/Y _08861_/X VGND VGND VPWR VPWR _08862_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08793_ _10013_/A _08793_/B VGND VGND VPWR VPWR _08793_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09414_ _09415_/A _09415_/B VGND VGND VPWR VPWR _09414_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09345_ _08703_/A _09791_/C _09937_/A _08509_/A VGND VGND VPWR VPWR _09345_/X sky130_fd_sc_hd__a22o_1
X_09276_ _08610_/A _09803_/A _09220_/A VGND VGND VPWR VPWR _09276_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10120_ _10120_/A _10120_/B VGND VGND VPWR VPWR _10120_/X sky130_fd_sc_hd__or2_1
X_10051_ _10024_/X _10050_/Y _10024_/X _10050_/Y VGND VGND VPWR VPWR _10077_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14790_ _14790_/A _14790_/B VGND VGND VPWR VPWR _14790_/X sky130_fd_sc_hd__and2_1
X_13810_ _13810_/A _13769_/X VGND VGND VPWR VPWR _13810_/X sky130_fd_sc_hd__or2b_1
XFILLER_113_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13741_ _13763_/A _13763_/B VGND VGND VPWR VPWR _13819_/A sky130_fd_sc_hd__and2_1
X_10953_ _11988_/A _10953_/B VGND VGND VPWR VPWR _10953_/X sky130_fd_sc_hd__and2_1
XFILLER_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16460_ _08229_/A _16460_/D VGND VGND VPWR VPWR _16460_/Q sky130_fd_sc_hd__dfxtp_1
X_13672_ _13620_/X _13671_/Y _13620_/X _13671_/Y VGND VGND VPWR VPWR _13691_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10884_ _09409_/A _09409_/B _09409_/Y VGND VGND VPWR VPWR _10885_/A sky130_fd_sc_hd__a21oi_1
X_16391_ _16389_/X _16390_/Y _16389_/X _16390_/Y VGND VGND VPWR VPWR _16392_/C sky130_fd_sc_hd__a2bb2o_1
X_12623_ _12623_/A _12623_/B VGND VGND VPWR VPWR _12623_/X sky130_fd_sc_hd__or2_1
X_15411_ _15450_/A _15409_/X _15410_/X VGND VGND VPWR VPWR _15411_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12554_ _12554_/A VGND VGND VPWR VPWR _12554_/Y sky130_fd_sc_hd__inv_2
X_15342_ _15375_/A _15340_/X _15341_/X VGND VGND VPWR VPWR _15342_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15273_ _15324_/A _15271_/X _15272_/X VGND VGND VPWR VPWR _15273_/Y sky130_fd_sc_hd__o21ai_1
X_11505_ _11504_/A _11504_/B _11504_/X _11303_/X VGND VGND VPWR VPWR _11632_/A sky130_fd_sc_hd__o22a_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14224_ _14090_/Y _14223_/X _14090_/Y _14223_/X VGND VGND VPWR VPWR _14225_/B sky130_fd_sc_hd__a2bb2oi_1
X_12485_ _14066_/A _12404_/B _12404_/Y _12356_/X VGND VGND VPWR VPWR _12485_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_8_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11436_ _13396_/A _11440_/B VGND VGND VPWR VPWR _11436_/Y sky130_fd_sc_hd__nor2_1
X_11367_ _12306_/A VGND VGND VPWR VPWR _14126_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14155_ _14153_/X _14154_/Y _14153_/X _14154_/Y VGND VGND VPWR VPWR _14155_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_125_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14086_ _14049_/X _14085_/X _14049_/X _14085_/X VGND VGND VPWR VPWR _14086_/Y sky130_fd_sc_hd__a2bb2oi_1
X_13106_ _13092_/Y _13104_/X _13105_/Y VGND VGND VPWR VPWR _13106_/X sky130_fd_sc_hd__o21a_1
X_10318_ _10299_/X _10317_/X _10299_/X _10317_/X VGND VGND VPWR VPWR _10319_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13037_ _14976_/A _13127_/B VGND VGND VPWR VPWR _13037_/Y sky130_fd_sc_hd__nor2_1
X_11298_ _11298_/A _11298_/B VGND VGND VPWR VPWR _11298_/Y sky130_fd_sc_hd__nor2_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10249_ _10247_/A _10247_/B _10247_/X _10248_/Y VGND VGND VPWR VPWR _10252_/B sky130_fd_sc_hd__o22ai_2
XFILLER_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14988_ _14979_/X _14987_/X _14979_/X _14987_/X VGND VGND VPWR VPWR _14988_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13939_ _15396_/A _13938_/B _13937_/X _13938_/X VGND VGND VPWR VPWR _13939_/X sky130_fd_sc_hd__o22a_1
X_15609_ _15609_/A VGND VGND VPWR VPWR _15609_/Y sky130_fd_sc_hd__inv_2
X_09130_ _09130_/A VGND VGND VPWR VPWR _09130_/Y sky130_fd_sc_hd__inv_2
X_09061_ _08823_/X _09044_/X _08823_/X _09044_/X VGND VGND VPWR VPWR _10017_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09963_ _09963_/A VGND VGND VPWR VPWR _09963_/Y sky130_fd_sc_hd__inv_2
X_08914_ _09066_/A VGND VGND VPWR VPWR _09401_/A sky130_fd_sc_hd__inv_2
XFILLER_131_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09884_/A _09884_/B _09885_/B VGND VGND VPWR VPWR _09908_/A sky130_fd_sc_hd__a21bo_1
XFILLER_85_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08944_/A _08719_/B _08719_/Y VGND VGND VPWR VPWR _09826_/B sky130_fd_sc_hd__a21oi_2
X_08776_ _08778_/B VGND VGND VPWR VPWR _08776_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09328_ _09328_/A _09328_/B VGND VGND VPWR VPWR _09328_/X sky130_fd_sc_hd__or2_1
X_09259_ _08904_/X _08809_/Y _10073_/A _09258_/X VGND VGND VPWR VPWR _09259_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12270_ _12270_/A VGND VGND VPWR VPWR _12270_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11221_ _12221_/A VGND VGND VPWR VPWR _14032_/A sky130_fd_sc_hd__buf_1
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11152_ _11152_/A VGND VGND VPWR VPWR _11152_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10103_ _10103_/A _10103_/B VGND VGND VPWR VPWR _10123_/B sky130_fd_sc_hd__nand2_1
XFILLER_122_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15960_ _15960_/A _15960_/B VGND VGND VPWR VPWR _15960_/X sky130_fd_sc_hd__or2_1
X_11083_ _13918_/A _11083_/B VGND VGND VPWR VPWR _11083_/X sky130_fd_sc_hd__or2_1
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15891_ _15877_/Y _15889_/X _15890_/Y VGND VGND VPWR VPWR _15891_/X sky130_fd_sc_hd__o21a_1
X_14911_ _14895_/Y _14909_/X _14910_/Y VGND VGND VPWR VPWR _14911_/X sky130_fd_sc_hd__o21a_1
X_10034_ _10034_/A _10034_/B VGND VGND VPWR VPWR _10034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14842_ _14841_/A _14841_/B _14841_/Y VGND VGND VPWR VPWR _14842_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14773_ _14742_/X _14772_/X _14742_/X _14772_/X VGND VGND VPWR VPWR _14774_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11985_ _11985_/A _11985_/B VGND VGND VPWR VPWR _11985_/X sky130_fd_sc_hd__or2_1
X_13724_ _13724_/A _13703_/X VGND VGND VPWR VPWR _13724_/X sky130_fd_sc_hd__or2b_1
X_10936_ _10936_/A VGND VGND VPWR VPWR _10936_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16443_ _16441_/Y _16442_/Y _16441_/Y _16442_/Y VGND VGND VPWR VPWR _16443_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10867_ _10867_/A _10867_/B VGND VGND VPWR VPWR _10867_/X sky130_fd_sc_hd__and2_1
X_13655_ _13703_/A _13703_/B VGND VGND VPWR VPWR _13724_/A sky130_fd_sc_hd__and2_1
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _11420_/X _12606_/B VGND VGND VPWR VPWR _12607_/B sky130_fd_sc_hd__and2b_1
XFILLER_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16374_ _16357_/X _16461_/Q _16358_/X _16397_/C _16361_/X VGND VGND VPWR VPWR _16461_/D
+ sky130_fd_sc_hd__o221a_2
X_13586_ _13581_/X _13585_/Y _13581_/X _13585_/Y VGND VGND VPWR VPWR _13642_/B sky130_fd_sc_hd__a2bb2o_1
X_10798_ _10798_/A _10798_/B VGND VGND VPWR VPWR _10798_/Y sky130_fd_sc_hd__nand2_1
X_12537_ _13438_/A _11384_/B _11384_/Y VGND VGND VPWR VPWR _12538_/B sky130_fd_sc_hd__o21a_1
X_15325_ _15271_/X _15324_/X _15271_/X _15324_/X VGND VGND VPWR VPWR _15331_/B sky130_fd_sc_hd__a2bb2o_1
X_15256_ _15202_/A _15202_/B _15202_/Y VGND VGND VPWR VPWR _15256_/Y sky130_fd_sc_hd__o21ai_1
X_12468_ _12437_/X _12467_/X _12437_/X _12467_/X VGND VGND VPWR VPWR _12468_/X sky130_fd_sc_hd__a2bb2o_1
X_14207_ _14207_/A _14207_/B VGND VGND VPWR VPWR _15869_/A sky130_fd_sc_hd__or2_1
X_11419_ _13405_/A _11420_/B VGND VGND VPWR VPWR _12606_/B sky130_fd_sc_hd__or2_1
XFILLER_99_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15187_ _15187_/A _15187_/B VGND VGND VPWR VPWR _15187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14138_ _14138_/A VGND VGND VPWR VPWR _14864_/A sky130_fd_sc_hd__inv_2
XFILLER_99_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12399_ _12359_/X _12398_/X _12359_/X _12398_/X VGND VGND VPWR VPWR _12401_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_98_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14069_ _14147_/A _14067_/X _14068_/X VGND VGND VPWR VPWR _14069_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08630_ _09225_/A VGND VGND VPWR VPWR _10017_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08561_ _08561_/A VGND VGND VPWR VPWR _08561_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08492_ _08321_/A _08251_/B _08472_/Y _08538_/A VGND VGND VPWR VPWR _08527_/A sky130_fd_sc_hd__o22a_1
XFILLER_35_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09113_ _09717_/A _09113_/B VGND VGND VPWR VPWR _09113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09044_ _08717_/A _08717_/B _08717_/X _09043_/Y VGND VGND VPWR VPWR _09044_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09946_ _09946_/A VGND VGND VPWR VPWR _09946_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09869_/X _08773_/Y _09869_/X _08773_/Y VGND VGND VPWR VPWR _09886_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08828_ _09458_/A VGND VGND VPWR VPWR _09500_/A sky130_fd_sc_hd__buf_1
X_08759_ _09331_/B VGND VGND VPWR VPWR _10133_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11770_ _11770_/A _11770_/B VGND VGND VPWR VPWR _11770_/X sky130_fd_sc_hd__and2_1
XFILLER_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10721_ _09975_/A _09650_/B _09650_/Y VGND VGND VPWR VPWR _10723_/A sky130_fd_sc_hd__o21ai_1
XFILLER_26_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13440_/A _13440_/B VGND VGND VPWR VPWR _13440_/Y sky130_fd_sc_hd__nand2_1
X_10652_ _10651_/Y _10534_/X _10579_/Y VGND VGND VPWR VPWR _10652_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13371_ _13371_/A _13371_/B VGND VGND VPWR VPWR _13371_/X sky130_fd_sc_hd__or2_1
X_10583_ _09723_/A _09723_/B _09723_/Y VGND VGND VPWR VPWR _10584_/A sky130_fd_sc_hd__o21ai_1
X_16090_ _16086_/Y _16223_/A _16089_/Y VGND VGND VPWR VPWR _16094_/B sky130_fd_sc_hd__o21ai_1
X_12322_ _12322_/A _12322_/B VGND VGND VPWR VPWR _12322_/X sky130_fd_sc_hd__and2_1
X_15110_ _15110_/A _15110_/B VGND VGND VPWR VPWR _15110_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12253_ _12252_/Y _12159_/X _12193_/Y VGND VGND VPWR VPWR _12253_/X sky130_fd_sc_hd__o21a_1
X_15041_ _15064_/A _15039_/X _15040_/X VGND VGND VPWR VPWR _15041_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11204_ _11204_/A _11089_/X VGND VGND VPWR VPWR _11204_/X sky130_fd_sc_hd__or2b_1
XFILLER_107_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12184_ _12261_/B _12183_/Y _12261_/B _12183_/Y VGND VGND VPWR VPWR _12259_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11135_ _12170_/A VGND VGND VPWR VPWR _13504_/A sky130_fd_sc_hd__buf_1
XFILLER_1_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15943_ _15886_/A _15886_/B _15886_/Y VGND VGND VPWR VPWR _15943_/Y sky130_fd_sc_hd__o21ai_1
X_11066_ _11244_/A VGND VGND VPWR VPWR _12232_/B sky130_fd_sc_hd__inv_2
XFILLER_95_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10017_ _10017_/A _10017_/B VGND VGND VPWR VPWR _10065_/B sky130_fd_sc_hd__nor2_1
X_15874_ _15892_/A _15892_/B VGND VGND VPWR VPWR _15874_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14825_ _14782_/A _14782_/B _14782_/X _14824_/X VGND VGND VPWR VPWR _14825_/X sky130_fd_sc_hd__o22a_1
XFILLER_91_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14756_ _14751_/X _14755_/X _14751_/X _14755_/X VGND VGND VPWR VPWR _14757_/B sky130_fd_sc_hd__a2bb2o_1
X_11968_ _11968_/A _11968_/B VGND VGND VPWR VPWR _11968_/Y sky130_fd_sc_hd__nand2_1
X_13707_ _13705_/Y _13706_/Y _13652_/Y VGND VGND VPWR VPWR _13778_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10919_ _14615_/A _10919_/B VGND VGND VPWR VPWR _10919_/X sky130_fd_sc_hd__or2_1
X_14687_ _15349_/A _14743_/B VGND VGND VPWR VPWR _14687_/Y sky130_fd_sc_hd__nand2_1
X_11899_ _11879_/Y _11897_/Y _11898_/Y VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__o21ai_1
X_16426_ _16426_/A _16434_/A VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__or2b_1
X_13638_ _15125_/A _13638_/B VGND VGND VPWR VPWR _13638_/Y sky130_fd_sc_hd__nand2_1
X_16357_ _16357_/A VGND VGND VPWR VPWR _16357_/X sky130_fd_sc_hd__buf_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13569_ _13569_/A VGND VGND VPWR VPWR _13569_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15308_ _15343_/A _15343_/B VGND VGND VPWR VPWR _15372_/A sky130_fd_sc_hd__and2_1
X_16288_ _16266_/A _16332_/A _16266_/Y VGND VGND VPWR VPWR _16288_/Y sky130_fd_sc_hd__o21ai_1
X_15239_ _15226_/X _15238_/Y _15226_/X _15238_/Y VGND VGND VPWR VPWR _15240_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09800_ _09800_/A _09834_/A VGND VGND VPWR VPWR _09801_/B sky130_fd_sc_hd__or2_1
XFILLER_101_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09731_ _09731_/A _09731_/B VGND VGND VPWR VPWR _09734_/B sky130_fd_sc_hd__or2_1
XFILLER_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09662_ _09993_/A _09662_/B VGND VGND VPWR VPWR _09662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08613_ _08612_/A _08354_/Y _08612_/Y _08354_/A VGND VGND VPWR VPWR _08614_/B sky130_fd_sc_hd__o22a_1
X_09593_ _09512_/X _09592_/X _09512_/X _09592_/X VGND VGND VPWR VPWR _09986_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _09860_/A VGND VGND VPWR VPWR _09740_/A sky130_fd_sc_hd__inv_2
XFILLER_63_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08475_ input15/X input31/X VGND VGND VPWR VPWR _08475_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09027_ _09005_/Y _08657_/Y _09005_/Y _08657_/Y VGND VGND VPWR VPWR _09028_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_123_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09929_ _09348_/B _09924_/Y _09863_/B VGND VGND VPWR VPWR _09929_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12940_ _12940_/A _12940_/B VGND VGND VPWR VPWR _12940_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12871_ _14757_/A _12944_/B VGND VGND VPWR VPWR _12871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14610_ _15347_/A _14662_/B VGND VGND VPWR VPWR _14610_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11822_ _11775_/A _11775_/B _11775_/A _11775_/B VGND VGND VPWR VPWR _11822_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15590_ _15590_/A _14394_/X VGND VGND VPWR VPWR _15590_/X sky130_fd_sc_hd__or2b_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14541_/A _14522_/X VGND VGND VPWR VPWR _14541_/X sky130_fd_sc_hd__or2b_1
X_11753_ _11772_/B VGND VGND VPWR VPWR _11753_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10704_ _11939_/A _10704_/B VGND VGND VPWR VPWR _10704_/Y sky130_fd_sc_hd__nand2_1
X_14472_ _15038_/A _11914_/Y _11862_/Y _14437_/X VGND VGND VPWR VPWR _14472_/X sky130_fd_sc_hd__o22a_1
X_11684_ _12428_/A _11623_/A _11624_/Y _11627_/X VGND VGND VPWR VPWR _11684_/X sky130_fd_sc_hd__o22a_1
X_16211_ _16255_/A _16322_/A VGND VGND VPWR VPWR _16211_/Y sky130_fd_sc_hd__nor2_1
X_13423_ _14101_/A _13426_/B VGND VGND VPWR VPWR _13423_/Y sky130_fd_sc_hd__nor2_1
X_10635_ _10735_/A _10635_/B VGND VGND VPWR VPWR _10635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16142_ _15712_/X _16142_/B VGND VGND VPWR VPWR _16142_/X sky130_fd_sc_hd__and2b_1
X_13354_ _15473_/A _13355_/B VGND VGND VPWR VPWR _13403_/A sky130_fd_sc_hd__and2_1
XFILLER_10_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12305_ _12245_/X _12304_/Y _12245_/X _12304_/Y VGND VGND VPWR VPWR _12306_/B sky130_fd_sc_hd__a2bb2o_1
X_10566_ _10566_/A VGND VGND VPWR VPWR _10566_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16073_ _16110_/A _16110_/B VGND VGND VPWR VPWR _16073_/X sky130_fd_sc_hd__and2_1
XFILLER_114_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13285_ _14731_/A _13285_/B VGND VGND VPWR VPWR _13285_/Y sky130_fd_sc_hd__nand2_1
X_10497_ _13621_/A _10529_/B VGND VGND VPWR VPWR _10497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12236_ _13351_/A _12236_/B VGND VGND VPWR VPWR _12236_/Y sky130_fd_sc_hd__nand2_1
X_15024_ _15030_/A _15030_/B VGND VGND VPWR VPWR _15079_/A sky130_fd_sc_hd__and2_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12167_ _12167_/A _12167_/B VGND VGND VPWR VPWR _12167_/X sky130_fd_sc_hd__or2_1
XFILLER_122_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11118_ _09782_/A _09782_/B _09782_/Y VGND VGND VPWR VPWR _11119_/A sky130_fd_sc_hd__o21ai_1
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12098_ _12160_/A _12160_/B VGND VGND VPWR VPWR _12098_/Y sky130_fd_sc_hd__nand2_1
X_15926_ _15897_/X _15925_/Y _15897_/X _15925_/Y VGND VGND VPWR VPWR _15960_/B sky130_fd_sc_hd__a2bb2o_1
Xinput7 wbs_adr_i[14] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_4
X_11049_ _15081_/A VGND VGND VPWR VPWR _14427_/A sky130_fd_sc_hd__buf_1
XFILLER_49_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15857_ _15857_/A VGND VGND VPWR VPWR _15902_/A sky130_fd_sc_hd__inv_2
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14808_ _14724_/X _14807_/X _14724_/X _14807_/X VGND VGND VPWR VPWR _14809_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15788_ _16089_/A _15788_/B VGND VGND VPWR VPWR _15788_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14739_ _14739_/A _14739_/B VGND VGND VPWR VPWR _14739_/X sky130_fd_sc_hd__or2_1
X_08260_ input15/X _08260_/B VGND VGND VPWR VPWR _08337_/A sky130_fd_sc_hd__nor2_1
X_16409_ _16409_/A VGND VGND VPWR VPWR _16409_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09714_ _09714_/A _09714_/B VGND VGND VPWR VPWR _09714_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09645_ _09960_/A _09645_/B VGND VGND VPWR VPWR _09645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09576_ _09515_/X _09575_/X _09515_/X _09575_/X VGND VGND VPWR VPWR _09995_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08527_/A VGND VGND VPWR VPWR _08527_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08458_ _08532_/B _08453_/Y _09331_/A VGND VGND VPWR VPWR _08459_/A sky130_fd_sc_hd__o21ai_1
XFILLER_11_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10420_ _10903_/A _10420_/B VGND VGND VPWR VPWR _12232_/A sky130_fd_sc_hd__nand2_2
X_08389_ _08389_/A VGND VGND VPWR VPWR _08389_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10351_ _10521_/A VGND VGND VPWR VPWR _10620_/A sky130_fd_sc_hd__inv_2
X_13070_ _13070_/A _13022_/X VGND VGND VPWR VPWR _13070_/X sky130_fd_sc_hd__or2b_1
X_10282_ _10282_/A VGND VGND VPWR VPWR _10282_/Y sky130_fd_sc_hd__inv_2
X_12021_ _11973_/X _12020_/Y _11973_/X _12020_/Y VGND VGND VPWR VPWR _12059_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13972_ _13972_/A VGND VGND VPWR VPWR _13973_/B sky130_fd_sc_hd__inv_2
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15711_ _15695_/X _15710_/Y _15695_/X _15710_/Y VGND VGND VPWR VPWR _15821_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12923_ _12923_/A VGND VGND VPWR VPWR _14459_/A sky130_fd_sc_hd__buf_1
XFILLER_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15642_ _15640_/A _15641_/A _15640_/Y _15641_/Y _15571_/A VGND VGND VPWR VPWR _16032_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_61_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12854_ _12854_/A _12854_/B VGND VGND VPWR VPWR _12854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15573_ _15491_/X _15573_/B VGND VGND VPWR VPWR _15573_/X sky130_fd_sc_hd__and2b_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12785_ _12785_/A _12785_/B VGND VGND VPWR VPWR _12785_/Y sky130_fd_sc_hd__nand2_1
X_11805_ _11805_/A _11805_/B VGND VGND VPWR VPWR _11805_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14524_/A VGND VGND VPWR VPWR _15190_/A sky130_fd_sc_hd__buf_1
X_11736_ _11742_/A _11743_/A VGND VGND VPWR VPWR _11736_/Y sky130_fd_sc_hd__nor2_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11667_ _12486_/A VGND VGND VPWR VPWR _15433_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14455_ _13274_/A _14429_/B _14429_/Y VGND VGND VPWR VPWR _14455_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14386_ _14386_/A _15956_/A VGND VGND VPWR VPWR _14386_/X sky130_fd_sc_hd__or2_1
X_13406_ _13406_/A _13406_/B VGND VGND VPWR VPWR _14240_/A sky130_fd_sc_hd__or2_2
X_10618_ _10618_/A _12605_/A VGND VGND VPWR VPWR _15212_/A sky130_fd_sc_hd__or2_1
X_11598_ _11574_/Y _10122_/Y _10237_/X VGND VGND VPWR VPWR _11599_/B sky130_fd_sc_hd__o21a_1
XFILLER_128_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16125_ _16125_/A _16125_/B VGND VGND VPWR VPWR _16386_/B sky130_fd_sc_hd__or2_1
X_13337_ _13337_/A _13337_/B VGND VGND VPWR VPWR _13337_/X sky130_fd_sc_hd__and2_1
X_10549_ _11850_/A VGND VGND VPWR VPWR _13516_/A sky130_fd_sc_hd__buf_1
X_16056_ _16059_/A _16054_/X _16055_/X VGND VGND VPWR VPWR _16056_/X sky130_fd_sc_hd__o21a_1
X_13268_ _13274_/A _13274_/B VGND VGND VPWR VPWR _13268_/Y sky130_fd_sc_hd__nor2_1
X_15007_ _12180_/X _15006_/X _12180_/X _15006_/X VGND VGND VPWR VPWR _15046_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12219_ _12219_/A _12143_/X VGND VGND VPWR VPWR _12219_/X sky130_fd_sc_hd__or2b_1
X_13199_ _13156_/Y _13197_/X _13198_/Y VGND VGND VPWR VPWR _13199_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15909_ _15856_/Y _15907_/X _15908_/Y VGND VGND VPWR VPWR _15909_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09430_ _09430_/A _09430_/B VGND VGND VPWR VPWR _09430_/X sky130_fd_sc_hd__or2_1
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09361_ _09478_/B _09863_/A _09347_/A VGND VGND VPWR VPWR _09361_/X sky130_fd_sc_hd__o21a_1
X_08312_ _08312_/A _08312_/B VGND VGND VPWR VPWR _08313_/A sky130_fd_sc_hd__or2_1
X_09292_ _08935_/A _08398_/Y _09235_/A _09628_/A VGND VGND VPWR VPWR _09293_/A sky130_fd_sc_hd__a31o_1
X_08243_ input5/X VGND VGND VPWR VPWR _08311_/A sky130_fd_sc_hd__inv_2
XFILLER_20_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09628_ _09628_/A _09628_/B VGND VGND VPWR VPWR _09628_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09559_ _08692_/A _09154_/A _09528_/Y _09558_/X VGND VGND VPWR VPWR _09559_/X sky130_fd_sc_hd__o22a_1
X_12570_ _14912_/A _12339_/B _12339_/Y VGND VGND VPWR VPWR _12571_/A sky130_fd_sc_hd__o21ai_1
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11521_ _10086_/X _11520_/X _10086_/X _11520_/X VGND VGND VPWR VPWR _11522_/B sky130_fd_sc_hd__a2bb2o_1
X_14240_ _14240_/A VGND VGND VPWR VPWR _14244_/B sky130_fd_sc_hd__inv_2
XFILLER_109_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11452_ _12349_/A VGND VGND VPWR VPWR _15540_/A sky130_fd_sc_hd__buf_1
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14171_ _14171_/A _12639_/X VGND VGND VPWR VPWR _14171_/X sky130_fd_sc_hd__or2b_1
X_11383_ _11257_/X _11382_/Y _11257_/X _11382_/Y VGND VGND VPWR VPWR _11384_/B sky130_fd_sc_hd__a2bb2o_1
X_10403_ _10403_/A VGND VGND VPWR VPWR _10403_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13122_ _13052_/Y _13120_/X _13121_/Y VGND VGND VPWR VPWR _13122_/X sky130_fd_sc_hd__o21a_1
X_10334_ _13530_/A VGND VGND VPWR VPWR _15028_/A sky130_fd_sc_hd__buf_1
XFILLER_127_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13053_ _13053_/A VGND VGND VPWR VPWR _13773_/A sky130_fd_sc_hd__inv_2
XFILLER_3_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _10197_/Y _10264_/Y _10197_/Y _10264_/Y VGND VGND VPWR VPWR _10265_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12004_ _11984_/X _12003_/X _11984_/X _12003_/X VGND VGND VPWR VPWR _12071_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10196_ _09342_/X _10195_/Y _09342_/X _10195_/Y VGND VGND VPWR VPWR _10196_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13955_ _13905_/Y _13953_/X _13954_/Y VGND VGND VPWR VPWR _13955_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13886_ _14832_/A _13991_/B VGND VGND VPWR VPWR _13886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12906_ _12839_/X _12905_/Y _12839_/X _12905_/Y VGND VGND VPWR VPWR _12926_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _15625_/A VGND VGND VPWR VPWR _15625_/Y sky130_fd_sc_hd__inv_2
X_12837_ _15087_/A _12836_/B _12835_/X _12836_/X VGND VGND VPWR VPWR _12837_/X sky130_fd_sc_hd__o22a_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _15556_/A _15556_/B VGND VGND VPWR VPWR _15556_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12768_ _12753_/Y _12766_/X _12767_/Y VGND VGND VPWR VPWR _12768_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15487_ _15434_/Y _15486_/X _15434_/Y _15486_/X VGND VGND VPWR VPWR _15554_/B sky130_fd_sc_hd__a2bb2o_1
X_14507_ _13002_/X _14506_/X _13002_/X _14506_/X VGND VGND VPWR VPWR _14508_/B sky130_fd_sc_hd__a2bb2o_1
X_11719_ _11719_/A _11719_/B VGND VGND VPWR VPWR _11719_/Y sky130_fd_sc_hd__nor2_1
X_12699_ _10310_/Y _12658_/Y _10310_/Y _12658_/Y VGND VGND VPWR VPWR _12700_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput21 wbs_dat_i[12] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_4
X_14438_ _11863_/Y _14437_/X _11863_/Y _14437_/X VGND VGND VPWR VPWR _14439_/B sky130_fd_sc_hd__o2bb2a_1
Xinput10 wbs_adr_i[2] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_4
Xinput32 wbs_dat_i[8] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__buf_4
X_14369_ _14376_/A _14376_/B VGND VGND VPWR VPWR _14370_/A sky130_fd_sc_hd__or2_1
X_16108_ _16108_/A _16108_/B VGND VGND VPWR VPWR _16179_/B sky130_fd_sc_hd__or2_1
XFILLER_116_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16039_ _16013_/Y _16037_/X _16038_/Y VGND VGND VPWR VPWR _16039_/X sky130_fd_sc_hd__o21a_1
XFILLER_103_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08930_ _08930_/A _10287_/A VGND VGND VPWR VPWR _08931_/A sky130_fd_sc_hd__or2_2
XFILLER_69_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08861_ _09496_/A _08817_/A _08819_/Y _08860_/X VGND VGND VPWR VPWR _08861_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08792_ _08793_/B VGND VGND VPWR VPWR _08792_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09413_ _09286_/Y _10876_/A _09412_/X VGND VGND VPWR VPWR _09415_/B sky130_fd_sc_hd__o21ai_1
XFILLER_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09344_ _09340_/X _09343_/X _09340_/X _09343_/X VGND VGND VPWR VPWR _09344_/X sky130_fd_sc_hd__o2bb2a_2
X_09275_ _09275_/A _09275_/B VGND VGND VPWR VPWR _09275_/X sky130_fd_sc_hd__or2_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10050_ _10050_/A _10050_/B VGND VGND VPWR VPWR _10050_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13740_ _13692_/X _13739_/X _13692_/X _13739_/X VGND VGND VPWR VPWR _13763_/B sky130_fd_sc_hd__a2bb2o_1
X_10952_ _10951_/A _10951_/B _10951_/X _10796_/X VGND VGND VPWR VPWR _10952_/X sky130_fd_sc_hd__o22a_1
XFILLER_43_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15410_ _15410_/A _15410_/B VGND VGND VPWR VPWR _15410_/X sky130_fd_sc_hd__or2_1
X_10883_ _10883_/A _10883_/B VGND VGND VPWR VPWR _10883_/X sky130_fd_sc_hd__and2_1
X_13671_ _15137_/A _13622_/B _13622_/Y VGND VGND VPWR VPWR _13671_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16390_ _16278_/A _16339_/X _16277_/X VGND VGND VPWR VPWR _16390_/Y sky130_fd_sc_hd__o21ai_1
X_12622_ _14220_/A _12620_/X _12621_/X VGND VGND VPWR VPWR _12622_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12553_ _12627_/A _12627_/B VGND VGND VPWR VPWR _14202_/A sky130_fd_sc_hd__and2_1
X_15341_ _15341_/A _15341_/B VGND VGND VPWR VPWR _15341_/X sky130_fd_sc_hd__or2_1
XFILLER_12_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15272_ _15272_/A _15272_/B VGND VGND VPWR VPWR _15272_/X sky130_fd_sc_hd__or2_1
X_11504_ _11504_/A _11504_/B VGND VGND VPWR VPWR _11504_/X sky130_fd_sc_hd__and2_1
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14223_ _14088_/X _14223_/B VGND VGND VPWR VPWR _14223_/X sky130_fd_sc_hd__and2b_1
X_12484_ _12486_/A _12486_/B VGND VGND VPWR VPWR _12484_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11435_ _11431_/Y _12574_/A _11434_/Y VGND VGND VPWR VPWR _11440_/B sky130_fd_sc_hd__o21ai_1
XFILLER_125_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11366_ _11569_/A _11366_/B VGND VGND VPWR VPWR _12306_/A sky130_fd_sc_hd__or2_1
X_14154_ _12426_/A _11615_/A _11616_/Y _13493_/X VGND VGND VPWR VPWR _14154_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_113_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14085_ _14812_/A _14043_/B _14043_/Y VGND VGND VPWR VPWR _14085_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13105_ _13747_/A _13105_/B VGND VGND VPWR VPWR _13105_/Y sky130_fd_sc_hd__nand2_1
X_10317_ _10367_/A _12700_/A _10316_/Y VGND VGND VPWR VPWR _10317_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11297_ _11297_/A VGND VGND VPWR VPWR _11297_/Y sky130_fd_sc_hd__inv_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13036_ _12952_/X _13035_/X _12952_/X _13035_/X VGND VGND VPWR VPWR _13127_/B sky130_fd_sc_hd__a2bb2o_1
X_10248_ _10248_/A VGND VGND VPWR VPWR _10248_/Y sky130_fd_sc_hd__inv_2
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10179_ _10180_/A _10180_/B VGND VGND VPWR VPWR _10179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14987_ _14981_/X _14986_/X _14981_/X _14986_/X VGND VGND VPWR VPWR _14987_/X sky130_fd_sc_hd__a2bb2o_1
X_13938_ _15396_/A _13938_/B VGND VGND VPWR VPWR _13938_/X sky130_fd_sc_hd__and2_1
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13869_ _11273_/A _13786_/B _13868_/Y _13783_/X VGND VGND VPWR VPWR _13869_/X sky130_fd_sc_hd__o22a_1
X_15608_ _14916_/A _15540_/B _15540_/Y VGND VGND VPWR VPWR _15609_/A sky130_fd_sc_hd__o21ai_1
X_15539_ _15539_/A VGND VGND VPWR VPWR _15539_/Y sky130_fd_sc_hd__inv_2
X_09060_ _08814_/X _09045_/X _08814_/X _09045_/X VGND VGND VPWR VPWR _10016_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09962_ _09962_/A VGND VGND VPWR VPWR _09962_/Y sky130_fd_sc_hd__inv_2
X_08913_ _09041_/A _08913_/B VGND VGND VPWR VPWR _09066_/A sky130_fd_sc_hd__or2_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09885_/A _09885_/B _09886_/B VGND VGND VPWR VPWR _09913_/A sky130_fd_sc_hd__a21bo_1
XFILLER_85_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08844_/A _10123_/A VGND VGND VPWR VPWR _08844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08775_ _10131_/A VGND VGND VPWR VPWR _08778_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09327_ _10241_/A VGND VGND VPWR VPWR _09328_/B sky130_fd_sc_hd__buf_1
XFILLER_21_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09258_ _08819_/A _08817_/A _10069_/A _09257_/X VGND VGND VPWR VPWR _09258_/X sky130_fd_sc_hd__o22a_1
X_09189_ _09189_/A VGND VGND VPWR VPWR _09190_/B sky130_fd_sc_hd__inv_2
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11220_ _13337_/A VGND VGND VPWR VPWR _12221_/A sky130_fd_sc_hd__inv_2
XFILLER_122_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11151_ _12268_/A _11314_/B _11150_/Y VGND VGND VPWR VPWR _11152_/A sky130_fd_sc_hd__o21ai_2
XFILLER_107_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10102_ _10102_/A _10102_/B VGND VGND VPWR VPWR _10103_/B sky130_fd_sc_hd__nor2_1
X_11082_ _11228_/A _11080_/X _11081_/X VGND VGND VPWR VPWR _11082_/X sky130_fd_sc_hd__o21a_1
X_14910_ _14910_/A _14910_/B VGND VGND VPWR VPWR _14910_/Y sky130_fd_sc_hd__nand2_1
X_15890_ _15890_/A _15890_/B VGND VGND VPWR VPWR _15890_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10033_ _09339_/X _10008_/X _10030_/Y _10032_/Y VGND VGND VPWR VPWR _10034_/B sky130_fd_sc_hd__a31o_1
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14841_ _14841_/A _14841_/B VGND VGND VPWR VPWR _14841_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14772_ _14772_/A _14771_/X VGND VGND VPWR VPWR _14772_/X sky130_fd_sc_hd__or2b_1
X_11984_ _13548_/A _11983_/B _11983_/X _11912_/X VGND VGND VPWR VPWR _11984_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13723_ _13775_/A _13775_/B VGND VGND VPWR VPWR _13801_/A sky130_fd_sc_hd__and2_1
X_10935_ _12068_/A _10935_/B VGND VGND VPWR VPWR _10935_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16442_ _16415_/X _16420_/X _16426_/X VGND VGND VPWR VPWR _16442_/Y sky130_fd_sc_hd__a21boi_1
X_10866_ _10773_/X _10865_/Y _10773_/X _10865_/Y VGND VGND VPWR VPWR _10867_/B sky130_fd_sc_hd__o2bb2a_1
X_13654_ _13705_/A _13653_/Y _13705_/A _13653_/Y VGND VGND VPWR VPWR _13703_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16373_ _16321_/X _16372_/Y _16321_/X _16372_/Y VGND VGND VPWR VPWR _16397_/C sky130_fd_sc_hd__a2bb2o_1
X_12605_ _12605_/A _12605_/B _13406_/B VGND VGND VPWR VPWR _14244_/A sky130_fd_sc_hd__and3_1
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15324_ _15324_/A _15272_/X VGND VGND VPWR VPWR _15324_/X sky130_fd_sc_hd__or2b_1
X_13585_ _13584_/A _13584_/B _13645_/A VGND VGND VPWR VPWR _13585_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10797_ _09263_/A _09263_/B _09263_/X VGND VGND VPWR VPWR _10798_/B sky130_fd_sc_hd__a21boi_1
X_12536_ _14114_/A VGND VGND VPWR VPWR _13438_/A sky130_fd_sc_hd__buf_1
XFILLER_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15255_ _15255_/A _15255_/B VGND VGND VPWR VPWR _15255_/Y sky130_fd_sc_hd__nand2_1
X_12467_ _12474_/A _12465_/X _12466_/X VGND VGND VPWR VPWR _12467_/X sky130_fd_sc_hd__o21a_1
X_14206_ _14105_/Y _14205_/X _14105_/Y _14205_/X VGND VGND VPWR VPWR _14207_/B sky130_fd_sc_hd__a2bb2oi_1
X_11418_ _11249_/X _11417_/X _11249_/X _11417_/X VGND VGND VPWR VPWR _11420_/B sky130_fd_sc_hd__a2bb2o_1
X_15186_ _15155_/X _15185_/Y _15155_/X _15185_/Y VGND VGND VPWR VPWR _15187_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14137_ _14138_/A _14139_/A VGND VGND VPWR VPWR _14137_/Y sky130_fd_sc_hd__nor2_1
X_12398_ _12398_/A _12397_/X VGND VGND VPWR VPWR _12398_/X sky130_fd_sc_hd__or2b_1
XFILLER_125_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11349_ _13890_/A _11350_/B VGND VGND VPWR VPWR _11351_/A sky130_fd_sc_hd__and2_1
XFILLER_4_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14068_ _14068_/A _14068_/B VGND VGND VPWR VPWR _14068_/X sky130_fd_sc_hd__or2_1
X_13019_ _13080_/A _13017_/X _13018_/X VGND VGND VPWR VPWR _13019_/X sky130_fd_sc_hd__o21a_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08560_ _08688_/A _10117_/B VGND VGND VPWR VPWR _08886_/A sky130_fd_sc_hd__nor2_1
X_08491_ _08326_/A _08254_/B _08473_/Y _08549_/A VGND VGND VPWR VPWR _08538_/A sky130_fd_sc_hd__o22a_1
XFILLER_90_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09112_ _09112_/A VGND VGND VPWR VPWR _09112_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09043_ _08718_/Y _09042_/X _08724_/X VGND VGND VPWR VPWR _09043_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09945_ _10252_/A _09310_/B _09310_/Y VGND VGND VPWR VPWR _09947_/A sky130_fd_sc_hd__o21ai_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09870_/X _08765_/Y _09870_/X _08765_/Y VGND VGND VPWR VPWR _09887_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _10017_/A _10125_/A VGND VGND VPWR VPWR _08827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08758_ _08757_/A _08745_/A _08757_/Y _08745_/Y VGND VGND VPWR VPWR _09331_/B sky130_fd_sc_hd__o22a_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08689_ _08886_/A _08687_/X _08886_/B VGND VGND VPWR VPWR _08689_/X sky130_fd_sc_hd__o21ba_1
XFILLER_26_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _11945_/A _10720_/B VGND VGND VPWR VPWR _10720_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10651_ _13633_/A _10651_/B VGND VGND VPWR VPWR _10651_/Y sky130_fd_sc_hd__nor2_1
X_13370_ _13382_/A _13368_/X _13369_/X VGND VGND VPWR VPWR _13370_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10582_ _11907_/A _10644_/B VGND VGND VPWR VPWR _10582_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12321_ _14082_/A _12318_/B _12319_/Y _12609_/A VGND VGND VPWR VPWR _12322_/B sky130_fd_sc_hd__o22a_1
X_12252_ _12252_/A _12252_/B VGND VGND VPWR VPWR _12252_/Y sky130_fd_sc_hd__nor2_1
X_15040_ _15040_/A _15040_/B VGND VGND VPWR VPWR _15040_/X sky130_fd_sc_hd__or2_1
X_11203_ _14056_/A VGND VGND VPWR VPWR _15452_/A sky130_fd_sc_hd__buf_1
XFILLER_79_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12183_ _12781_/A _12262_/A _12182_/Y VGND VGND VPWR VPWR _12183_/Y sky130_fd_sc_hd__a21oi_1
X_11134_ _10083_/A _11133_/Y _09966_/Y _11133_/A _10957_/X VGND VGND VPWR VPWR _12170_/A
+ sky130_fd_sc_hd__o221a_1
X_15942_ _15950_/A _15950_/B VGND VGND VPWR VPWR _16020_/A sky130_fd_sc_hd__and2_1
X_11065_ _11065_/A _11065_/B VGND VGND VPWR VPWR _11244_/A sky130_fd_sc_hd__or2_1
XFILLER_95_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10016_ _10016_/A _10016_/B VGND VGND VPWR VPWR _10069_/B sky130_fd_sc_hd__nor2_1
X_15873_ _14214_/X _15843_/X _14214_/X _15843_/X VGND VGND VPWR VPWR _15892_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14824_ _14786_/A _14786_/B _14786_/X _14823_/X VGND VGND VPWR VPWR _14824_/X sky130_fd_sc_hd__o22a_1
XFILLER_63_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11967_ _11954_/Y _11965_/X _11966_/Y VGND VGND VPWR VPWR _11967_/X sky130_fd_sc_hd__o21a_1
X_14755_ _14754_/A _14754_/B _14754_/Y VGND VGND VPWR VPWR _14755_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10918_ _10918_/A VGND VGND VPWR VPWR _14615_/A sky130_fd_sc_hd__buf_1
X_13706_ _13706_/A _13706_/B VGND VGND VPWR VPWR _13706_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16425_ _16416_/Y _16437_/B _16415_/A VGND VGND VPWR VPWR _16434_/A sky130_fd_sc_hd__a21oi_1
X_14686_ _14666_/X _14685_/Y _14666_/X _14685_/Y VGND VGND VPWR VPWR _14743_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11898_ _12990_/A _11898_/B VGND VGND VPWR VPWR _11898_/Y sky130_fd_sc_hd__nand2_1
X_10849_ _12061_/A VGND VGND VPWR VPWR _10918_/A sky130_fd_sc_hd__inv_2
X_13637_ _13637_/A VGND VGND VPWR VPWR _15125_/A sky130_fd_sc_hd__buf_1
X_16356_ _08230_/X _16466_/Q _08233_/X _16402_/B _16343_/X VGND VGND VPWR VPWR _16466_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_118_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13568_ _13568_/A _13568_/B VGND VGND VPWR VPWR _13569_/A sky130_fd_sc_hd__nand2_1
X_16287_ _16334_/A _16334_/B VGND VGND VPWR VPWR _16287_/Y sky130_fd_sc_hd__nor2_1
X_12519_ _12635_/A _12635_/B VGND VGND VPWR VPWR _14178_/A sky130_fd_sc_hd__and2_1
X_15307_ _15278_/X _15306_/Y _15278_/X _15306_/Y VGND VGND VPWR VPWR _15343_/B sky130_fd_sc_hd__a2bb2o_1
X_15238_ _15184_/A _15184_/B _15184_/Y VGND VGND VPWR VPWR _15238_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13499_ _13501_/A VGND VGND VPWR VPWR _15051_/A sky130_fd_sc_hd__buf_1
XFILLER_8_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15169_ _15107_/A _15107_/B _15107_/Y _15099_/X VGND VGND VPWR VPWR _15169_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09730_ _09730_/A _09730_/B VGND VGND VPWR VPWR _09733_/A sky130_fd_sc_hd__or2_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09661_ _09591_/Y _09659_/X _09660_/Y VGND VGND VPWR VPWR _09661_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08612_ _08612_/A VGND VGND VPWR VPWR _08612_/Y sky130_fd_sc_hd__inv_2
X_09592_ _09490_/A _09490_/B _09490_/Y VGND VGND VPWR VPWR _09592_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08543_ _08543_/A _08543_/B VGND VGND VPWR VPWR _09860_/A sky130_fd_sc_hd__or2_2
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08474_ input16/X input32/X VGND VGND VPWR VPWR _08474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09026_ _08645_/X _09007_/Y _08645_/X _09007_/Y VGND VGND VPWR VPWR _09539_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09928_ _09928_/A _09928_/B VGND VGND VPWR VPWR _09931_/A sky130_fd_sc_hd__and2_1
XFILLER_105_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09859_ _09859_/A _09859_/B VGND VGND VPWR VPWR _09914_/A sky130_fd_sc_hd__or2_1
XFILLER_105_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12870_ _12857_/X _12869_/Y _12857_/X _12869_/Y VGND VGND VPWR VPWR _12944_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11821_ _13625_/A _11841_/B VGND VGND VPWR VPWR _11821_/Y sky130_fd_sc_hd__nor2_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _15249_/A VGND VGND VPWR VPWR _14586_/A sky130_fd_sc_hd__buf_1
XFILLER_121_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11752_ _11757_/B _11751_/X _11757_/B _11751_/X VGND VGND VPWR VPWR _11772_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14439_/A _14439_/B _14436_/X _14439_/Y VGND VGND VPWR VPWR _14471_/X sky130_fd_sc_hd__o2bb2a_1
X_10703_ _10782_/A _10702_/Y _10782_/A _10702_/Y VGND VGND VPWR VPWR _10704_/B sky130_fd_sc_hd__a2bb2o_1
X_11683_ _15163_/A VGND VGND VPWR VPWR _12428_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16210_ _16255_/B VGND VGND VPWR VPWR _16322_/A sky130_fd_sc_hd__buf_1
X_13422_ _13418_/Y _13420_/Y _13421_/Y VGND VGND VPWR VPWR _13426_/B sky130_fd_sc_hd__o21ai_2
X_10634_ _10634_/A VGND VGND VPWR VPWR _10634_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16141_ _16140_/A _16139_/Y _16140_/Y _16139_/A _16388_/A VGND VGND VPWR VPWR _16273_/A
+ sky130_fd_sc_hd__a221o_1
X_13353_ _11413_/X _13352_/X _11413_/X _13352_/X VGND VGND VPWR VPWR _13355_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12304_ _14015_/A _12206_/B _12206_/Y VGND VGND VPWR VPWR _12304_/Y sky130_fd_sc_hd__o21ai_1
X_10565_ _11920_/A _10673_/B _10564_/Y VGND VGND VPWR VPWR _10566_/A sky130_fd_sc_hd__o21ai_2
X_16072_ _16041_/X _16071_/Y _16041_/X _16071_/Y VGND VGND VPWR VPWR _16110_/B sky130_fd_sc_hd__a2bb2o_1
X_13284_ _13284_/A VGND VGND VPWR VPWR _13284_/Y sky130_fd_sc_hd__inv_2
X_10496_ _10434_/X _10495_/X _10434_/X _10495_/X VGND VGND VPWR VPWR _10529_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12235_ _12235_/A VGND VGND VPWR VPWR _12235_/X sky130_fd_sc_hd__buf_1
XFILLER_107_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15023_ _11737_/Y _14998_/X _11737_/Y _14998_/X VGND VGND VPWR VPWR _15030_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12166_ _13649_/A _12165_/B _12165_/X _12074_/X VGND VGND VPWR VPWR _12166_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11117_ _11115_/Y _11116_/Y _10995_/Y VGND VGND VPWR VPWR _11289_/A sky130_fd_sc_hd__o21ai_1
X_12097_ _12072_/X _12096_/Y _12072_/X _12096_/Y VGND VGND VPWR VPWR _12160_/B sky130_fd_sc_hd__a2bb2o_1
X_15925_ _15898_/A _15898_/B _15898_/Y VGND VGND VPWR VPWR _15925_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11048_ _12840_/A VGND VGND VPWR VPWR _15081_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 wbs_adr_i[15] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__buf_1
X_15856_ _15908_/A _15908_/B VGND VGND VPWR VPWR _15856_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14807_ _14807_/A _14807_/B VGND VGND VPWR VPWR _14807_/X sky130_fd_sc_hd__or2_1
XFILLER_91_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15787_ _15787_/A VGND VGND VPWR VPWR _16089_/A sky130_fd_sc_hd__buf_1
X_12999_ _12922_/A _12998_/Y _12922_/A _12998_/Y VGND VGND VPWR VPWR _13010_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14738_ _14784_/A _14736_/X _14737_/X VGND VGND VPWR VPWR _14738_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14669_ _14669_/A VGND VGND VPWR VPWR _15184_/A sky130_fd_sc_hd__buf_1
XFILLER_32_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16408_ _16399_/Y _16407_/Y _16393_/Y VGND VGND VPWR VPWR _16409_/A sky130_fd_sc_hd__o21ai_1
X_16339_ _16281_/Y _16337_/X _16338_/Y VGND VGND VPWR VPWR _16339_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09713_ _09713_/A VGND VGND VPWR VPWR _09714_/B sky130_fd_sc_hd__inv_2
XFILLER_95_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09644_ _09544_/X _09643_/X _09544_/X _09643_/X VGND VGND VPWR VPWR _10731_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ _09484_/A _09484_/B _09484_/Y VGND VGND VPWR VPWR _09575_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08526_ _08694_/A _10120_/B VGND VGND VPWR VPWR _08871_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08457_ _10009_/A VGND VGND VPWR VPWR _09331_/A sky130_fd_sc_hd__inv_2
XFILLER_51_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08388_ _08388_/A VGND VGND VPWR VPWR _08388_/Y sky130_fd_sc_hd__inv_2
X_10350_ _10350_/A _10350_/B VGND VGND VPWR VPWR _10521_/A sky130_fd_sc_hd__or2_1
XFILLER_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10281_ _10281_/A VGND VGND VPWR VPWR _10350_/A sky130_fd_sc_hd__inv_2
XFILLER_3_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09009_ _08962_/X _09025_/S _08631_/Y VGND VGND VPWR VPWR _09024_/S sky130_fd_sc_hd__o21ai_1
X_12020_ _13068_/A _11974_/B _11974_/Y VGND VGND VPWR VPWR _12020_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13971_ _13969_/X _13970_/Y _13969_/X _13970_/Y VGND VGND VPWR VPWR _13972_/A sky130_fd_sc_hd__a2bb2o_1
X_15710_ _16055_/A _15696_/B _15696_/Y VGND VGND VPWR VPWR _15710_/Y sky130_fd_sc_hd__o21ai_1
X_12922_ _12922_/A VGND VGND VPWR VPWR _12922_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15641_ _15641_/A VGND VGND VPWR VPWR _15641_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12853_ _12804_/Y _12851_/X _12852_/Y VGND VGND VPWR VPWR _12853_/X sky130_fd_sc_hd__o21a_1
X_15572_ _15595_/A VGND VGND VPWR VPWR _15700_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12729_/Y _12782_/X _12783_/Y VGND VGND VPWR VPWR _12784_/X sky130_fd_sc_hd__o21a_1
X_11804_ _11803_/A _11803_/B _11803_/X _11764_/B VGND VGND VPWR VPWR _11852_/B sky130_fd_sc_hd__a22o_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14541_/A _14521_/X _14522_/X VGND VGND VPWR VPWR _14523_/X sky130_fd_sc_hd__o21a_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11735_ _10226_/X _11745_/B _10226_/A _11745_/B VGND VGND VPWR VPWR _11743_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _14461_/A _14461_/B VGND VGND VPWR VPWR _14454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13405_ _13405_/A _13405_/B VGND VGND VPWR VPWR _13405_/X sky130_fd_sc_hd__and2_1
X_11666_ _09199_/Y _11663_/Y _09199_/A _11663_/A _11665_/X VGND VGND VPWR VPWR _12486_/A
+ sky130_fd_sc_hd__a221o_4
X_14385_ _15628_/A _14383_/X _14384_/X VGND VGND VPWR VPWR _14385_/X sky130_fd_sc_hd__o21a_1
X_10617_ _10522_/A _10616_/Y _10522_/A _10616_/Y VGND VGND VPWR VPWR _10626_/B sky130_fd_sc_hd__a2bb2o_1
X_11597_ _15163_/A VGND VGND VPWR VPWR _12410_/A sky130_fd_sc_hd__inv_2
X_16124_ _16061_/X _16122_/X _16133_/B VGND VGND VPWR VPWR _16124_/X sky130_fd_sc_hd__o21a_1
X_13336_ _13281_/A _13335_/Y _13281_/A _13335_/Y VGND VGND VPWR VPWR _13337_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10548_ _09700_/A _10547_/Y _09700_/Y _10547_/A _10957_/A VGND VGND VPWR VPWR _11850_/A
+ sky130_fd_sc_hd__o221a_1
X_16055_ _16055_/A _16055_/B VGND VGND VPWR VPWR _16055_/X sky130_fd_sc_hd__or2_1
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13267_ _13183_/X _13266_/Y _13183_/X _13266_/Y VGND VGND VPWR VPWR _13274_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12218_ _12218_/A _12218_/B VGND VGND VPWR VPWR _12218_/Y sky130_fd_sc_hd__nand2_1
X_10479_ _10443_/X _10478_/X _10443_/X _10478_/X VGND VGND VPWR VPWR _10538_/B sky130_fd_sc_hd__a2bb2o_1
X_15006_ _12088_/A _15005_/X _12087_/X VGND VGND VPWR VPWR _15006_/X sky130_fd_sc_hd__o21a_1
X_13198_ _13198_/A _13198_/B VGND VGND VPWR VPWR _13198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12149_ _13906_/A _12149_/B VGND VGND VPWR VPWR _12149_/X sky130_fd_sc_hd__or2_1
XFILLER_69_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15908_ _15908_/A _15908_/B VGND VGND VPWR VPWR _15908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15839_ _15839_/A _15839_/B VGND VGND VPWR VPWR _15840_/A sky130_fd_sc_hd__or2_1
XFILLER_92_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09360_ _09345_/X _09359_/X _09345_/X _09359_/X VGND VGND VPWR VPWR _09360_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08311_ _08311_/A input21/X VGND VGND VPWR VPWR _08312_/B sky130_fd_sc_hd__nor2_1
X_09291_ _10230_/A VGND VGND VPWR VPWR _09298_/A sky130_fd_sc_hd__buf_1
XFILLER_60_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08242_ _08242_/A input6/X VGND VGND VPWR VPWR _08307_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09627_ _09627_/A VGND VGND VPWR VPWR _09707_/A sky130_fd_sc_hd__inv_2
XFILLER_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09558_ _08690_/A _09017_/A _09530_/Y _09557_/X VGND VGND VPWR VPWR _09558_/X sky130_fd_sc_hd__o22a_1
XFILLER_70_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08509_ _08509_/A VGND VGND VPWR VPWR _08656_/A sky130_fd_sc_hd__inv_2
XFILLER_24_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11520_ _10037_/X _11520_/B VGND VGND VPWR VPWR _11520_/X sky130_fd_sc_hd__and2b_1
X_09489_ _08789_/A _09469_/X _08789_/A _09469_/X VGND VGND VPWR VPWR _09490_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11451_ _11256_/X _11450_/Y _11256_/X _11450_/Y VGND VGND VPWR VPWR _12544_/A sky130_fd_sc_hd__a2bb2o_1
X_14170_ _14282_/A _14170_/B VGND VGND VPWR VPWR _15910_/A sky130_fd_sc_hd__or2_1
XFILLER_109_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11382_ _14056_/A _11206_/B _11206_/Y VGND VGND VPWR VPWR _11382_/Y sky130_fd_sc_hd__o21ai_1
X_10402_ _10402_/A VGND VGND VPWR VPWR _10402_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13121_ _15240_/A _13121_/B VGND VGND VPWR VPWR _13121_/Y sky130_fd_sc_hd__nand2_1
X_10333_ _11783_/A VGND VGND VPWR VPWR _13530_/A sky130_fd_sc_hd__buf_1
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13052_ _15240_/A _13121_/B VGND VGND VPWR VPWR _13052_/Y sky130_fd_sc_hd__nor2_1
X_10264_ _11574_/A _10237_/B _10237_/X _11599_/A VGND VGND VPWR VPWR _10264_/Y sky130_fd_sc_hd__a22oi_1
X_12003_ _11007_/A _12073_/B _11007_/A _12073_/B VGND VGND VPWR VPWR _12003_/X sky130_fd_sc_hd__a2bb2o_1
X_10195_ _10122_/Y _10193_/Y _10194_/Y VGND VGND VPWR VPWR _10195_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13954_ _15412_/A _13954_/B VGND VGND VPWR VPWR _13954_/Y sky130_fd_sc_hd__nand2_1
X_13885_ _13862_/X _13884_/X _13862_/X _13884_/X VGND VGND VPWR VPWR _13991_/B sky130_fd_sc_hd__a2bb2o_1
X_12905_ _12840_/A _12840_/B _12840_/Y VGND VGND VPWR VPWR _12905_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _15624_/A VGND VGND VPWR VPWR _15624_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12836_ _12836_/A _12836_/B VGND VGND VPWR VPWR _12836_/X sky130_fd_sc_hd__and2_1
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15488_/Y _15553_/Y _15554_/Y VGND VGND VPWR VPWR _15555_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _13610_/Y _13616_/A _15146_/A _13616_/Y VGND VGND VPWR VPWR _14506_/X sky130_fd_sc_hd__a22o_1
X_12767_ _12767_/A _12767_/B VGND VGND VPWR VPWR _12767_/Y sky130_fd_sc_hd__nand2_1
X_15486_ _14930_/A _15437_/B _15437_/X _15485_/X VGND VGND VPWR VPWR _15486_/X sky130_fd_sc_hd__o22a_1
X_11718_ _12831_/A _11716_/A _10425_/A _11717_/Y VGND VGND VPWR VPWR _11719_/B sky130_fd_sc_hd__o22a_1
X_12698_ _12698_/A _12698_/B VGND VGND VPWR VPWR _12698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput11 wbs_adr_i[3] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_4
X_11649_ _12393_/A _11649_/B VGND VGND VPWR VPWR _11649_/Y sky130_fd_sc_hd__nor2_1
X_14437_ _15036_/A _11848_/Y _11813_/Y _14419_/X VGND VGND VPWR VPWR _14437_/X sky130_fd_sc_hd__o22a_1
Xinput22 wbs_dat_i[13] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_2
X_14368_ _14368_/A _14368_/B VGND VGND VPWR VPWR _14376_/B sky130_fd_sc_hd__nor2_1
Xinput33 wbs_dat_i[9] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_4
X_16107_ _16079_/X _16105_/X _16187_/B VGND VGND VPWR VPWR _16107_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13319_ _13369_/A _13369_/B VGND VGND VPWR VPWR _13382_/A sky130_fd_sc_hd__and2_1
XFILLER_6_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14299_ _13445_/X _14298_/X _13445_/X _14298_/X VGND VGND VPWR VPWR _14300_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16038_ _16038_/A _16038_/B VGND VGND VPWR VPWR _16038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08860_ _09498_/A _08825_/A _08827_/Y _08859_/X VGND VGND VPWR VPWR _08860_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08791_ _10129_/A VGND VGND VPWR VPWR _08793_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09412_ _09412_/A _09412_/B VGND VGND VPWR VPWR _09412_/X sky130_fd_sc_hd__or2_1
XFILLER_80_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09343_ _09146_/X _09342_/B _09146_/X _09342_/X VGND VGND VPWR VPWR _09343_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09274_ _10244_/A VGND VGND VPWR VPWR _09275_/B sky130_fd_sc_hd__buf_1
XFILLER_33_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08989_ _08989_/A VGND VGND VPWR VPWR _08989_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10951_ _10951_/A _10951_/B VGND VGND VPWR VPWR _10951_/X sky130_fd_sc_hd__and2_1
XFILLER_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13670_ _13693_/A _13693_/B VGND VGND VPWR VPWR _13739_/A sky130_fd_sc_hd__and2_1
XFILLER_44_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12621_ _12621_/A _12621_/B VGND VGND VPWR VPWR _12621_/X sky130_fd_sc_hd__or2_1
X_10882_ _10771_/X _10881_/Y _10771_/X _10881_/Y VGND VGND VPWR VPWR _10883_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12552_ _12549_/Y _12551_/Y _12549_/A _12551_/A _12501_/A VGND VGND VPWR VPWR _12627_/B
+ sky130_fd_sc_hd__o221a_1
X_15340_ _15378_/A _15338_/X _15339_/X VGND VGND VPWR VPWR _15340_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12483_ _12477_/Y _12482_/Y _12477_/Y _12482_/Y VGND VGND VPWR VPWR _12486_/B sky130_fd_sc_hd__a2bb2o_1
X_15271_ _15270_/A _15270_/B _11064_/B _15270_/X VGND VGND VPWR VPWR _15271_/X sky130_fd_sc_hd__o22a_1
X_11503_ _12387_/A VGND VGND VPWR VPWR _13975_/A sky130_fd_sc_hd__buf_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14222_ _15875_/A _14257_/B VGND VGND VPWR VPWR _14222_/Y sky130_fd_sc_hd__nor2_1
X_11434_ _12575_/A _11434_/B VGND VGND VPWR VPWR _11434_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14153_ _14076_/Y _14152_/X _14076_/Y _14152_/X VGND VGND VPWR VPWR _14153_/X sky130_fd_sc_hd__a2bb2o_1
X_11365_ _08977_/X _11364_/X _08977_/X _11364_/X VGND VGND VPWR VPWR _11366_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_125_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14084_ _14084_/A _14084_/B VGND VGND VPWR VPWR _14084_/X sky130_fd_sc_hd__and2_1
X_13104_ _13095_/Y _13102_/X _13103_/Y VGND VGND VPWR VPWR _13104_/X sky130_fd_sc_hd__o21a_1
X_11296_ _11295_/Y _11123_/X _11164_/Y VGND VGND VPWR VPWR _11296_/X sky130_fd_sc_hd__o21a_1
X_10316_ _10367_/A _11757_/A VGND VGND VPWR VPWR _10316_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13035_ _13039_/A _13033_/X _13034_/X VGND VGND VPWR VPWR _13035_/X sky130_fd_sc_hd__o21a_1
X_10247_ _10247_/A _10247_/B VGND VGND VPWR VPWR _10247_/X sky130_fd_sc_hd__and2_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10178_ _10108_/A _10177_/Y _10106_/Y VGND VGND VPWR VPWR _10180_/B sky130_fd_sc_hd__o21ai_1
X_14986_ _14983_/Y _14985_/X _14983_/Y _14985_/X VGND VGND VPWR VPWR _14986_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13937_ _13937_/A VGND VGND VPWR VPWR _13937_/X sky130_fd_sc_hd__buf_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13868_ _13868_/A VGND VGND VPWR VPWR _13868_/Y sky130_fd_sc_hd__inv_2
X_15607_ _15679_/A _15679_/B VGND VGND VPWR VPWR _15607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13799_ _13776_/X _13798_/X _13776_/X _13798_/X VGND VGND VPWR VPWR _13860_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12819_ _12842_/A _12842_/B VGND VGND VPWR VPWR _12819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15538_ _15479_/Y _15537_/X _15479_/Y _15537_/X VGND VGND VPWR VPWR _15539_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15469_ _15397_/X _15468_/X _15397_/X _15468_/X VGND VGND VPWR VPWR _15470_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09961_ _09960_/A _09972_/B _09960_/Y VGND VGND VPWR VPWR _09962_/A sky130_fd_sc_hd__o21ai_1
X_08912_ _08970_/A _08970_/B VGND VGND VPWR VPWR _08912_/X sky130_fd_sc_hd__and2_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _09886_/A _09886_/B _09887_/B VGND VGND VPWR VPWR _09918_/A sky130_fd_sc_hd__a21bo_1
XFILLER_111_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _08843_/A VGND VGND VPWR VPWR _08844_/A sky130_fd_sc_hd__buf_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08774_ _08773_/A _08739_/A _08773_/Y _08739_/Y VGND VGND VPWR VPWR _10131_/A sky130_fd_sc_hd__o22a_1
XFILLER_85_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09326_ _09325_/X _08888_/Y _09325_/X _08888_/Y VGND VGND VPWR VPWR _10241_/A sky130_fd_sc_hd__o2bb2a_1
X_09257_ _08962_/X _08825_/A _10065_/A _09256_/X VGND VGND VPWR VPWR _09257_/X sky130_fd_sc_hd__o22a_1
X_09188_ _09561_/B _09156_/X _09561_/B _09156_/X VGND VGND VPWR VPWR _09189_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11150_ _12268_/A _11314_/B VGND VGND VPWR VPWR _11150_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10101_ _10099_/A _08679_/B _10100_/Y VGND VGND VPWR VPWR _10108_/A sky130_fd_sc_hd__a21oi_2
X_11081_ _13922_/A _11081_/B VGND VGND VPWR VPWR _11081_/X sky130_fd_sc_hd__or2_1
XFILLER_88_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10032_ _09339_/X _10008_/X _10030_/Y VGND VGND VPWR VPWR _10032_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14840_ _12383_/Y _14839_/X _12383_/Y _14839_/X VGND VGND VPWR VPWR _14841_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_90_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14771_ _14771_/A _14771_/B VGND VGND VPWR VPWR _14771_/X sky130_fd_sc_hd__or2_1
XFILLER_76_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13722_ _13704_/X _13721_/X _13704_/X _13721_/X VGND VGND VPWR VPWR _13775_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11983_ _13548_/A _11983_/B VGND VGND VPWR VPWR _11983_/X sky130_fd_sc_hd__and2_1
X_10934_ _12158_/A VGND VGND VPWR VPWR _13053_/A sky130_fd_sc_hd__buf_1
XFILLER_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16441_ _16416_/Y _16429_/B _16440_/X VGND VGND VPWR VPWR _16441_/Y sky130_fd_sc_hd__o21ai_1
X_10865_ _13073_/A _10720_/B _10720_/Y VGND VGND VPWR VPWR _10865_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13653_ _15119_/A _13706_/B _13652_/Y VGND VGND VPWR VPWR _13653_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _16322_/A _16322_/B _16322_/Y VGND VGND VPWR VPWR _16372_/Y sky130_fd_sc_hd__o21ai_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12604_ _12617_/A _12617_/B VGND VGND VPWR VPWR _12604_/X sky130_fd_sc_hd__and2_1
X_13584_ _13584_/A _13584_/B VGND VGND VPWR VPWR _13645_/A sky130_fd_sc_hd__nand2_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ _12631_/A _12631_/B VGND VGND VPWR VPWR _14190_/A sky130_fd_sc_hd__and2_1
X_15323_ _15333_/A _15333_/B VGND VGND VPWR VPWR _15387_/A sky130_fd_sc_hd__and2_1
X_10796_ _10795_/A _10795_/B _10795_/X _10658_/X VGND VGND VPWR VPWR _10796_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12466_ _13989_/A _12466_/B VGND VGND VPWR VPWR _12466_/X sky130_fd_sc_hd__or2_1
X_15254_ _15221_/X _15253_/Y _15221_/X _15253_/Y VGND VGND VPWR VPWR _15255_/B sky130_fd_sc_hd__a2bb2o_1
X_14205_ _14106_/A _14106_/B _14106_/Y VGND VGND VPWR VPWR _14205_/X sky130_fd_sc_hd__o21a_1
X_11417_ _11248_/X _11417_/B VGND VGND VPWR VPWR _11417_/X sky130_fd_sc_hd__and2b_1
X_12397_ _12397_/A _12397_/B VGND VGND VPWR VPWR _12397_/X sky130_fd_sc_hd__or2_1
X_15185_ _15119_/A _15119_/B _15119_/Y VGND VGND VPWR VPWR _15185_/Y sky130_fd_sc_hd__o21ai_1
X_14136_ _14063_/X _14135_/X _14063_/X _14135_/X VGND VGND VPWR VPWR _14139_/A sky130_fd_sc_hd__a2bb2o_1
X_11348_ _11277_/X _11347_/X _11277_/X _11347_/X VGND VGND VPWR VPWR _11350_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14067_ _14141_/A _14065_/X _14066_/X VGND VGND VPWR VPWR _14067_/X sky130_fd_sc_hd__o21a_1
X_11279_ _09438_/X _11278_/X _09438_/X _11278_/X VGND VGND VPWR VPWR _11280_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13018_ _14489_/A _13018_/B VGND VGND VPWR VPWR _13018_/X sky130_fd_sc_hd__or2_1
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14969_ _14929_/X _14968_/X _14929_/X _14968_/X VGND VGND VPWR VPWR _14996_/A sky130_fd_sc_hd__a2bb2oi_1
XFILLER_47_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08490_ _08331_/A _08257_/B _08474_/Y _08561_/A VGND VGND VPWR VPWR _08549_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09111_ _09538_/B _09031_/B _09032_/B VGND VGND VPWR VPWR _09112_/A sky130_fd_sc_hd__a21bo_1
XFILLER_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09042_ _08843_/A _09459_/B _08719_/Y _09064_/A VGND VGND VPWR VPWR _09042_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09944_ _11843_/A VGND VGND VPWR VPWR _13629_/A sky130_fd_sc_hd__buf_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _09871_/X _08757_/Y _09871_/X _08757_/Y VGND VGND VPWR VPWR _09888_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _09252_/B VGND VGND VPWR VPWR _10125_/A sky130_fd_sc_hd__buf_1
XFILLER_85_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08757_ _08757_/A VGND VGND VPWR VPWR _08757_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08688_ _08688_/A _10117_/B VGND VGND VPWR VPWR _08886_/B sky130_fd_sc_hd__and2_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10650_ _11867_/A VGND VGND VPWR VPWR _13633_/A sky130_fd_sc_hd__buf_1
XFILLER_110_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09309_ _10252_/A _09310_/B VGND VGND VPWR VPWR _09309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10581_ _10534_/X _10580_/Y _10534_/X _10580_/Y VGND VGND VPWR VPWR _10644_/B sky130_fd_sc_hd__a2bb2o_1
X_12320_ _12320_/A _13406_/B VGND VGND VPWR VPWR _12609_/A sky130_fd_sc_hd__or2_1
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12251_ _12290_/A VGND VGND VPWR VPWR _13204_/A sky130_fd_sc_hd__buf_1
XFILLER_79_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11202_ _14021_/A VGND VGND VPWR VPWR _14056_/A sky130_fd_sc_hd__buf_1
XFILLER_122_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12182_ _12781_/A _12262_/A VGND VGND VPWR VPWR _12182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11133_ _11133_/A VGND VGND VPWR VPWR _11133_/Y sky130_fd_sc_hd__inv_2
X_15941_ _15887_/X _15940_/Y _15887_/X _15940_/Y VGND VGND VPWR VPWR _15950_/B sky130_fd_sc_hd__a2bb2o_1
X_11064_ _12041_/B _11064_/B _13096_/A VGND VGND VPWR VPWR _11065_/B sky130_fd_sc_hd__and3_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10015_ _10015_/A _10015_/B VGND VGND VPWR VPWR _10073_/B sky130_fd_sc_hd__nor2_1
X_15872_ _15872_/A VGND VGND VPWR VPWR _15892_/A sky130_fd_sc_hd__inv_2
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14823_ _14790_/A _14790_/B _14790_/X _14822_/X VGND VGND VPWR VPWR _14823_/X sky130_fd_sc_hd__o22a_1
XFILLER_91_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11966_ _11966_/A _11966_/B VGND VGND VPWR VPWR _11966_/Y sky130_fd_sc_hd__nand2_1
X_14754_ _14754_/A _14754_/B VGND VGND VPWR VPWR _14754_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10917_ _11025_/A _10914_/X _10916_/X VGND VGND VPWR VPWR _10917_/X sky130_fd_sc_hd__o21a_1
X_14685_ _14746_/A _14746_/B _14684_/Y VGND VGND VPWR VPWR _14685_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13705_ _13705_/A VGND VGND VPWR VPWR _13705_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16424_ _16421_/Y _16447_/B _16447_/A _16415_/A _16420_/X VGND VGND VPWR VPWR _16426_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11897_ _11897_/A VGND VGND VPWR VPWR _11897_/Y sky130_fd_sc_hd__inv_2
X_13636_ _13636_/A VGND VGND VPWR VPWR _13636_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10848_ _09266_/A _10847_/A _09269_/A _10847_/Y _10926_/A VGND VGND VPWR VPWR _12061_/A
+ sky130_fd_sc_hd__a221o_2
X_16355_ _16331_/X _16354_/Y _16331_/X _16354_/Y VGND VGND VPWR VPWR _16402_/B sky130_fd_sc_hd__a2bb2o_1
X_13567_ _13532_/X _13566_/Y _13532_/X _13566_/Y VGND VGND VPWR VPWR _13568_/B sky130_fd_sc_hd__a2bb2o_1
X_10779_ _10930_/A _10779_/B VGND VGND VPWR VPWR _12066_/A sky130_fd_sc_hd__or2_2
XFILLER_12_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16286_ _16267_/X _16285_/Y _16267_/X _16285_/Y VGND VGND VPWR VPWR _16334_/B sky130_fd_sc_hd__o2bb2a_1
X_12518_ _12517_/A _12517_/B _12517_/Y _12501_/X VGND VGND VPWR VPWR _12635_/B sky130_fd_sc_hd__o211a_1
X_15306_ _14586_/A _15249_/B _15249_/Y VGND VGND VPWR VPWR _15306_/Y sky130_fd_sc_hd__o21ai_1
X_13498_ _15104_/A _13498_/B VGND VGND VPWR VPWR _13498_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15237_ _15237_/A _15237_/B VGND VGND VPWR VPWR _15237_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12449_ _13975_/A _12449_/B VGND VGND VPWR VPWR _12449_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15168_ _15167_/A _15167_/B _15167_/Y VGND VGND VPWR VPWR _15168_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14119_ _14120_/A _14121_/A VGND VGND VPWR VPWR _14119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15099_ _15054_/A _15054_/B _15054_/Y _15098_/X VGND VGND VPWR VPWR _15099_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09660_ _09990_/A _09660_/B VGND VGND VPWR VPWR _09660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08611_ _08611_/A VGND VGND VPWR VPWR _08611_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09591_ _09990_/A _09660_/B VGND VGND VPWR VPWR _09591_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08542_ _09472_/B VGND VGND VPWR VPWR _08690_/A sky130_fd_sc_hd__buf_1
XFILLER_35_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08473_ input17/X input33/X VGND VGND VPWR VPWR _08473_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09025_ _08632_/X _08962_/X _09025_/S VGND VGND VPWR VPWR _09538_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09927_ _11298_/B _09926_/X VGND VGND VPWR VPWR _09928_/B sky130_fd_sc_hd__or2b_1
XFILLER_131_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09858_ _09858_/A _09904_/A VGND VGND VPWR VPWR _09859_/B sky130_fd_sc_hd__or2_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09789_ _09753_/Y _11494_/A _09788_/X VGND VGND VPWR VPWR _09789_/X sky130_fd_sc_hd__o21a_1
X_08809_ _08810_/B VGND VGND VPWR VPWR _08809_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11820_ _11796_/X _11819_/X _11796_/X _11819_/X VGND VGND VPWR VPWR _11841_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11751_ _11751_/A _11750_/X VGND VGND VPWR VPWR _11751_/X sky130_fd_sc_hd__or2b_1
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10702_ _13699_/A _10781_/B _10701_/Y VGND VGND VPWR VPWR _10702_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11680_/Y _11681_/Y _11680_/Y _11681_/Y VGND VGND VPWR VPWR _11682_/X sky130_fd_sc_hd__o2bb2a_1
X_14470_ _14442_/Y _14468_/X _14469_/Y VGND VGND VPWR VPWR _14470_/X sky130_fd_sc_hd__o21a_1
X_13421_ _14096_/A _13421_/B VGND VGND VPWR VPWR _13421_/Y sky130_fd_sc_hd__nand2_1
X_10633_ _10606_/Y _10631_/Y _10632_/Y VGND VGND VPWR VPWR _10634_/A sky130_fd_sc_hd__o21ai_1
XFILLER_14_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16140_ _16140_/A VGND VGND VPWR VPWR _16140_/Y sky130_fd_sc_hd__inv_2
X_13352_ _14722_/A _13272_/B _13272_/Y VGND VGND VPWR VPWR _13352_/X sky130_fd_sc_hd__a21o_1
X_10564_ _11920_/A _10673_/B VGND VGND VPWR VPWR _10564_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16071_ _16042_/A _16042_/B _16042_/Y VGND VGND VPWR VPWR _16071_/Y sky130_fd_sc_hd__o21ai_1
X_12303_ _12303_/A _12303_/B VGND VGND VPWR VPWR _12303_/Y sky130_fd_sc_hd__nand2_1
X_13283_ _13255_/Y _13281_/Y _13282_/Y VGND VGND VPWR VPWR _13284_/A sky130_fd_sc_hd__o21ai_1
X_10495_ _10396_/A _10400_/B _10396_/A _10400_/B VGND VGND VPWR VPWR _10495_/X sky130_fd_sc_hd__a2bb2o_1
X_15022_ _15032_/A _15032_/B VGND VGND VPWR VPWR _15076_/A sky130_fd_sc_hd__and2_1
XFILLER_123_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12234_ _12232_/Y _12233_/X _12232_/Y _12233_/X VGND VGND VPWR VPWR _12236_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12165_ _13649_/A _12165_/B VGND VGND VPWR VPWR _12165_/X sky130_fd_sc_hd__and2_1
XFILLER_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11116_ _11116_/A VGND VGND VPWR VPWR _11116_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12096_ _13706_/A _12163_/B _12095_/Y VGND VGND VPWR VPWR _12096_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15924_ _15962_/A _15962_/B VGND VGND VPWR VPWR _16002_/A sky130_fd_sc_hd__and2_1
XFILLER_77_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11047_ _13568_/A VGND VGND VPWR VPWR _12840_/A sky130_fd_sc_hd__buf_1
X_15855_ _14284_/X _15850_/X _14284_/X _15850_/X VGND VGND VPWR VPWR _15908_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 wbs_adr_i[1] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_4
X_14806_ _14806_/A _14806_/B VGND VGND VPWR VPWR _14806_/X sky130_fd_sc_hd__and2_1
XFILLER_36_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15786_ _15666_/X _15785_/X _15666_/X _15785_/X VGND VGND VPWR VPWR _15786_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12998_ _14459_/A _12924_/B _12924_/Y VGND VGND VPWR VPWR _12998_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14737_ _14737_/A _14737_/B VGND VGND VPWR VPWR _14737_/X sky130_fd_sc_hd__or2_1
X_11949_ _12990_/A _11898_/B _11898_/Y VGND VGND VPWR VPWR _11949_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14668_ _14591_/X _14605_/A _14604_/X VGND VGND VPWR VPWR _14668_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16407_ _16407_/A _16407_/B _16407_/C _16407_/D VGND VGND VPWR VPWR _16407_/Y sky130_fd_sc_hd__nor4_1
X_13619_ _12923_/A _13609_/B _13609_/X _13618_/X VGND VGND VPWR VPWR _13619_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16338_ _16338_/A _16338_/B VGND VGND VPWR VPWR _16338_/Y sky130_fd_sc_hd__nand2_1
X_14599_ _14594_/X _14598_/X _14594_/X _14598_/X VGND VGND VPWR VPWR _14600_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16269_ _16162_/Y _16267_/X _16268_/Y VGND VGND VPWR VPWR _16269_/X sky130_fd_sc_hd__o21a_1
XFILLER_114_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09712_ _09686_/A _09686_/B _09689_/A VGND VGND VPWR VPWR _10216_/A sky130_fd_sc_hd__a21bo_1
XFILLER_68_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09643_ _09538_/A _09538_/B _09538_/X VGND VGND VPWR VPWR _09643_/X sky130_fd_sc_hd__o21ba_1
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09574_ _09997_/A _09666_/B VGND VGND VPWR VPWR _09574_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _08524_/A _08459_/Y _08524_/Y _08459_/A VGND VGND VPWR VPWR _10120_/B sky130_fd_sc_hd__o22a_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08456_ _08532_/A VGND VGND VPWR VPWR _10009_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08387_ _08387_/A _08387_/B VGND VGND VPWR VPWR _08388_/A sky130_fd_sc_hd__or2_1
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10280_ _11720_/A VGND VGND VPWR VPWR _13479_/A sky130_fd_sc_hd__buf_1
XFILLER_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09008_ _09500_/A _09228_/B _09007_/Y VGND VGND VPWR VPWR _09025_/S sky130_fd_sc_hd__o21ai_1
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13970_ _13874_/A _13869_/X _13874_/B VGND VGND VPWR VPWR _13970_/Y sky130_fd_sc_hd__o21bai_1
X_12921_ _13003_/A _12920_/B _13002_/A _12920_/Y VGND VGND VPWR VPWR _12922_/A sky130_fd_sc_hd__o2bb2a_1
X_15640_ _15640_/A VGND VGND VPWR VPWR _15640_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12852_ _12852_/A _12852_/B VGND VGND VPWR VPWR _12852_/Y sky130_fd_sc_hd__nand2_1
X_15571_ _15571_/A VGND VGND VPWR VPWR _15595_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12783_ _12783_/A _12783_/B VGND VGND VPWR VPWR _12783_/Y sky130_fd_sc_hd__nand2_1
X_11803_ _11803_/A _11803_/B VGND VGND VPWR VPWR _11803_/X sky130_fd_sc_hd__or2_1
XFILLER_42_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _15193_/A _14522_/B VGND VGND VPWR VPWR _14522_/X sky130_fd_sc_hd__or2_1
XFILLER_42_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11734_ _11733_/A _11733_/B _10213_/B _11733_/X VGND VGND VPWR VPWR _11745_/B sky130_fd_sc_hd__a22o_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14453_ _14432_/X _14452_/X _14432_/X _14452_/X VGND VGND VPWR VPWR _14461_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11665_ _11664_/A _11664_/B _09189_/A _09190_/B _11664_/Y VGND VGND VPWR VPWR _11665_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13404_ _13350_/Y _13403_/X _13350_/Y _13403_/X VGND VGND VPWR VPWR _13405_/B sky130_fd_sc_hd__a2bb2o_1
X_10616_ _11833_/A _10523_/B _10523_/Y VGND VGND VPWR VPWR _10616_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14384_ _14384_/A _15954_/A VGND VGND VPWR VPWR _14384_/X sky130_fd_sc_hd__or2_1
X_11596_ _09750_/B _11595_/Y _09749_/X _11595_/A _10957_/X VGND VGND VPWR VPWR _15163_/A
+ sky130_fd_sc_hd__o221a_1
X_16123_ _16123_/A _16123_/B VGND VGND VPWR VPWR _16133_/B sky130_fd_sc_hd__or2_1
X_13335_ _14729_/A _13282_/B _13282_/Y VGND VGND VPWR VPWR _13335_/Y sky130_fd_sc_hd__o21ai_1
X_10547_ _10547_/A VGND VGND VPWR VPWR _10547_/Y sky130_fd_sc_hd__inv_2
X_16054_ _15998_/X _16052_/Y _16062_/B VGND VGND VPWR VPWR _16054_/X sky130_fd_sc_hd__o21a_1
X_13266_ _15331_/A _13184_/B _13184_/Y VGND VGND VPWR VPWR _13266_/Y sky130_fd_sc_hd__o21ai_1
X_10478_ _13519_/A _10544_/B _13519_/A _10544_/B VGND VGND VPWR VPWR _10478_/X sky130_fd_sc_hd__a2bb2o_1
X_12217_ _12144_/X _12216_/X _12144_/X _12216_/X VGND VGND VPWR VPWR _12218_/B sky130_fd_sc_hd__a2bb2o_1
X_15005_ _11998_/A _15004_/X _11997_/X VGND VGND VPWR VPWR _15005_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13197_ _13159_/Y _13195_/X _13196_/Y VGND VGND VPWR VPWR _13197_/X sky130_fd_sc_hd__o21a_1
X_12148_ _12213_/A _12146_/X _12147_/X VGND VGND VPWR VPWR _12148_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12079_ _12167_/A VGND VGND VPWR VPWR _12779_/A sky130_fd_sc_hd__buf_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15907_ _15904_/Y _15905_/X _15906_/Y VGND VGND VPWR VPWR _15907_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15838_ _15838_/A VGND VGND VPWR VPWR _15839_/B sky130_fd_sc_hd__inv_2
XFILLER_18_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15769_ _14904_/A _14904_/B _14904_/Y VGND VGND VPWR VPWR _15770_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08310_ _08308_/Y _08309_/A _08308_/A _08309_/Y _08304_/X VGND VGND VPWR VPWR _08521_/B
+ sky130_fd_sc_hd__o221a_1
X_09290_ _08922_/B _08936_/Y _08922_/B _08936_/Y VGND VGND VPWR VPWR _10230_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08241_ input22/X VGND VGND VPWR VPWR _08242_/A sky130_fd_sc_hd__inv_2
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09626_ _08922_/A _09625_/Y _08922_/A _09625_/Y VGND VGND VPWR VPWR _09952_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_70_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09557_ _08688_/A _09019_/A _09532_/Y _09556_/X VGND VGND VPWR VPWR _09557_/X sky130_fd_sc_hd__o22a_1
X_09488_ _09488_/A _09488_/B VGND VGND VPWR VPWR _09488_/Y sky130_fd_sc_hd__nor2_1
X_08508_ _08508_/A VGND VGND VPWR VPWR _09346_/B sky130_fd_sc_hd__inv_2
XFILLER_24_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08439_ _08439_/A VGND VGND VPWR VPWR _08439_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11450_ _14109_/A _11212_/B _11212_/Y VGND VGND VPWR VPWR _11450_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11381_ _12312_/A VGND VGND VPWR VPWR _14114_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10401_ _09304_/A _10235_/A _09304_/Y VGND VGND VPWR VPWR _10403_/A sky130_fd_sc_hd__o21ai_1
X_13120_ _13057_/Y _13118_/X _13119_/Y VGND VGND VPWR VPWR _13120_/X sky130_fd_sc_hd__o21a_1
X_10332_ _11719_/A VGND VGND VPWR VPWR _11783_/A sky130_fd_sc_hd__buf_1
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13051_ _13029_/X _13050_/X _13029_/X _13050_/X VGND VGND VPWR VPWR _13121_/B sky130_fd_sc_hd__a2bb2o_1
X_12002_ _12075_/B _12001_/Y _12075_/B _12001_/Y VGND VGND VPWR VPWR _12073_/B sky130_fd_sc_hd__o2bb2a_1
X_10263_ _09371_/B _10238_/B _10238_/X _11533_/A VGND VGND VPWR VPWR _11599_/A sky130_fd_sc_hd__a22o_1
XFILLER_87_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10194_ _10194_/A _10194_/B VGND VGND VPWR VPWR _10194_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13953_ _13909_/Y _13951_/X _13952_/Y VGND VGND VPWR VPWR _13953_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13884_ _13884_/A _13883_/X VGND VGND VPWR VPWR _13884_/X sky130_fd_sc_hd__or2b_1
X_12904_ _12926_/A VGND VGND VPWR VPWR _14461_/A sky130_fd_sc_hd__buf_1
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _14912_/A _15529_/B _15529_/Y VGND VGND VPWR VPWR _15625_/A sky130_fd_sc_hd__o21ai_1
X_12835_ _12916_/A VGND VGND VPWR VPWR _12835_/X sky130_fd_sc_hd__buf_1
XFILLER_62_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15554_/A _15554_/B VGND VGND VPWR VPWR _15554_/Y sky130_fd_sc_hd__nand2_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14505_/A VGND VGND VPWR VPWR _15216_/A sky130_fd_sc_hd__buf_1
X_12766_ _12756_/Y _12764_/X _12765_/Y VGND VGND VPWR VPWR _12766_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15485_ _14774_/A _15440_/B _15440_/X _15484_/X VGND VGND VPWR VPWR _15485_/X sky130_fd_sc_hd__o22a_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11788_/A _11717_/B VGND VGND VPWR VPWR _11717_/Y sky130_fd_sc_hd__nor2_1
X_12697_ _10381_/A _12660_/A _10381_/Y _12660_/Y VGND VGND VPWR VPWR _12698_/B sky130_fd_sc_hd__o22a_1
Xinput12 wbs_adr_i[4] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_4
X_11648_ _11648_/A _11647_/X VGND VGND VPWR VPWR _11648_/X sky130_fd_sc_hd__or2b_1
X_14436_ _14421_/A _14421_/B _14421_/Y _14435_/X VGND VGND VPWR VPWR _14436_/X sky130_fd_sc_hd__o2bb2a_1
X_14367_ _14240_/A _14366_/A _14244_/B _14366_/Y VGND VGND VPWR VPWR _14368_/B sky130_fd_sc_hd__o22a_1
Xinput23 wbs_dat_i[14] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_4
X_11579_ _13133_/A VGND VGND VPWR VPWR _12788_/A sky130_fd_sc_hd__clkbuf_2
X_16106_ _16106_/A _16106_/B VGND VGND VPWR VPWR _16187_/B sky130_fd_sc_hd__or2_1
X_13318_ _13299_/A _13317_/Y _13299_/A _13317_/Y VGND VGND VPWR VPWR _13369_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14298_ _13446_/A _13446_/B _13446_/Y VGND VGND VPWR VPWR _14298_/X sky130_fd_sc_hd__o21a_1
X_16037_ _16016_/Y _16035_/X _16036_/Y VGND VGND VPWR VPWR _16037_/X sky130_fd_sc_hd__o21a_1
X_13249_ _13191_/X _13248_/Y _13191_/X _13248_/Y VGND VGND VPWR VPWR _13285_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08790_ _08789_/A _08733_/A _08789_/Y _08733_/Y VGND VGND VPWR VPWR _10129_/A sky130_fd_sc_hd__o22a_1
XFILLER_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09411_ _09412_/A _09412_/B VGND VGND VPWR VPWR _10876_/A sky130_fd_sc_hd__and2_1
X_09342_ _09342_/A _09342_/B VGND VGND VPWR VPWR _09342_/X sky130_fd_sc_hd__and2_1
XFILLER_21_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09273_ _09258_/X _08905_/Y _09258_/X _08905_/Y VGND VGND VPWR VPWR _10244_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08988_ _08468_/Y _08987_/X _08468_/Y _08987_/X VGND VGND VPWR VPWR _08988_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10950_ _12095_/A VGND VGND VPWR VPWR _13706_/A sky130_fd_sc_hd__buf_1
XFILLER_56_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10881_ _13083_/A _10738_/B _10738_/Y VGND VGND VPWR VPWR _10881_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09609_ _09981_/A _09654_/B VGND VGND VPWR VPWR _09609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12620_ _14226_/A _12618_/X _12619_/X VGND VGND VPWR VPWR _12620_/X sky130_fd_sc_hd__o21a_1
XFILLER_73_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12551_ _12551_/A VGND VGND VPWR VPWR _12551_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12482_ _13995_/A _12478_/B _12478_/Y VGND VGND VPWR VPWR _12482_/Y sky130_fd_sc_hd__o21ai_1
X_15270_ _15270_/A _15270_/B VGND VGND VPWR VPWR _15270_/X sky130_fd_sc_hd__and2_1
X_11502_ _12946_/A VGND VGND VPWR VPWR _12387_/A sky130_fd_sc_hd__inv_2
XFILLER_12_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14221_ _12620_/X _14220_/X _12620_/X _14220_/X VGND VGND VPWR VPWR _14257_/B sky130_fd_sc_hd__a2bb2o_1
X_11433_ _11253_/X _11432_/Y _11253_/X _11432_/Y VGND VGND VPWR VPWR _12574_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14152_ _14150_/X _14151_/X _14150_/X _14151_/X VGND VGND VPWR VPWR _14152_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11364_ _08890_/X _11364_/B VGND VGND VPWR VPWR _11364_/X sky130_fd_sc_hd__and2b_1
X_14083_ _14082_/A _14082_/B _14240_/A _14082_/Y VGND VGND VPWR VPWR _14084_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13103_ _14564_/A _13103_/B VGND VGND VPWR VPWR _13103_/Y sky130_fd_sc_hd__nand2_1
X_11295_ _12187_/A _11295_/B VGND VGND VPWR VPWR _11295_/Y sky130_fd_sc_hd__nor2_1
X_10315_ _11757_/A VGND VGND VPWR VPWR _12700_/A sky130_fd_sc_hd__buf_1
XFILLER_112_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13034_ _14836_/A _13034_/B VGND VGND VPWR VPWR _13034_/X sky130_fd_sc_hd__or2_1
X_10246_ _10235_/X _10175_/A _10234_/A VGND VGND VPWR VPWR _10247_/B sky130_fd_sc_hd__o21ai_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10177_ _10177_/A _10177_/B VGND VGND VPWR VPWR _10177_/Y sky130_fd_sc_hd__nor2_1
X_14985_ _14929_/X _14984_/Y _14967_/Y VGND VGND VPWR VPWR _14985_/X sky130_fd_sc_hd__o21a_1
X_13936_ _13936_/A _13936_/B VGND VGND VPWR VPWR _13937_/A sky130_fd_sc_hd__or2_1
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15606_ _14389_/X _15605_/X _14389_/X _15605_/X VGND VGND VPWR VPWR _15679_/B sky130_fd_sc_hd__a2bb2o_1
X_13867_ _13975_/A VGND VGND VPWR VPWR _15110_/A sky130_fd_sc_hd__buf_1
X_13798_ _13798_/A _13797_/X VGND VGND VPWR VPWR _13798_/X sky130_fd_sc_hd__or2b_1
XFILLER_62_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12818_ _12766_/X _12817_/Y _12766_/X _12817_/Y VGND VGND VPWR VPWR _12842_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15537_ _15455_/A _15455_/B _15455_/A _15455_/B VGND VGND VPWR VPWR _15537_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12711_/X _12748_/X _12711_/X _12748_/X VGND VGND VPWR VPWR _12769_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15468_ _15468_/A _15398_/X VGND VGND VPWR VPWR _15468_/X sky130_fd_sc_hd__or2b_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14419_ _15034_/A _11799_/Y _11767_/Y _14418_/X VGND VGND VPWR VPWR _14419_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15399_ _15468_/A _15397_/X _15398_/X VGND VGND VPWR VPWR _15399_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09960_ _09960_/A _09972_/B VGND VGND VPWR VPWR _09960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08911_ _08910_/Y _08860_/X _08910_/Y _08860_/X VGND VGND VPWR VPWR _08970_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09887_/A _09887_/B _09888_/B VGND VGND VPWR VPWR _09923_/A sky130_fd_sc_hd__a21bo_1
XFILLER_97_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _10123_/A VGND VGND VPWR VPWR _08842_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08773_/A VGND VGND VPWR VPWR _08773_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09325_ _08893_/X _08792_/Y _10047_/A _09260_/X VGND VGND VPWR VPWR _09325_/X sky130_fd_sc_hd__o22a_1
X_09256_ _10018_/A _08834_/A _10061_/A _09255_/Y VGND VGND VPWR VPWR _09256_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09187_ _09429_/A _09191_/B VGND VGND VPWR VPWR _11664_/A sky130_fd_sc_hd__nor2_1
XFILLER_107_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11080_ _11234_/A _11077_/X _11079_/X VGND VGND VPWR VPWR _11080_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10100_ _10110_/A VGND VGND VPWR VPWR _10100_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10031_ _10008_/A _10008_/B _10008_/X _10030_/Y VGND VGND VPWR VPWR _10031_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14770_ _14771_/A _14771_/B VGND VGND VPWR VPWR _14772_/A sky130_fd_sc_hd__and2_1
XFILLER_17_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13721_ _13721_/A _13720_/X VGND VGND VPWR VPWR _13721_/X sky130_fd_sc_hd__or2b_1
X_11982_ _11981_/Y _11910_/X _11933_/Y VGND VGND VPWR VPWR _11982_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10933_ _11587_/A _10933_/B VGND VGND VPWR VPWR _12158_/A sky130_fd_sc_hd__or2_1
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16440_ _16412_/Y _16415_/X _16437_/B _16447_/B VGND VGND VPWR VPWR _16440_/X sky130_fd_sc_hd__o22a_1
X_10864_ _10867_/A VGND VGND VPWR VPWR _14623_/A sky130_fd_sc_hd__buf_1
XFILLER_71_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13652_ _15119_/A _13706_/B VGND VGND VPWR VPWR _13652_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16371_ _16357_/X _16462_/Q _16358_/X _16397_/D _16361_/X VGND VGND VPWR VPWR _16462_/D
+ sky130_fd_sc_hd__o221a_2
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12603_ _12600_/Y _12602_/A _12600_/A _12602_/Y _12500_/A VGND VGND VPWR VPWR _12617_/B
+ sky130_fd_sc_hd__o221a_1
X_10795_ _10795_/A _10795_/B VGND VGND VPWR VPWR _10795_/X sky130_fd_sc_hd__and2_1
X_13583_ _13538_/X _13582_/Y _13538_/X _13582_/Y VGND VGND VPWR VPWR _13584_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _12533_/A _12533_/B _12533_/Y _12501_/X VGND VGND VPWR VPWR _12631_/B sky130_fd_sc_hd__o211a_1
X_15322_ _15273_/Y _15321_/X _15273_/Y _15321_/X VGND VGND VPWR VPWR _15333_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_40_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12465_ _12398_/A _12359_/X _12397_/X VGND VGND VPWR VPWR _12465_/X sky130_fd_sc_hd__o21a_1
X_15253_ _15199_/A _15199_/B _15199_/Y VGND VGND VPWR VPWR _15253_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14204_ _15866_/A _14266_/B VGND VGND VPWR VPWR _14204_/Y sky130_fd_sc_hd__nor2_1
X_12396_ _12397_/A _12397_/B VGND VGND VPWR VPWR _12398_/A sky130_fd_sc_hd__and2_1
X_15184_ _15184_/A _15184_/B VGND VGND VPWR VPWR _15184_/Y sky130_fd_sc_hd__nand2_1
X_11416_ _09403_/X _08931_/A _08931_/Y _10515_/Y _08997_/A VGND VGND VPWR VPWR _13405_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14135_ _14135_/A _14064_/X VGND VGND VPWR VPWR _14135_/X sky130_fd_sc_hd__or2b_1
X_11347_ _14745_/A _11480_/B _11480_/A _11480_/B VGND VGND VPWR VPWR _11347_/X sky130_fd_sc_hd__a2bb2o_1
X_14066_ _14066_/A _14066_/B VGND VGND VPWR VPWR _14066_/X sky130_fd_sc_hd__or2_1
XFILLER_79_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11278_ _09785_/A _09374_/A _09431_/X VGND VGND VPWR VPWR _11278_/X sky130_fd_sc_hd__o21a_1
X_13017_ _13085_/A _13014_/X _13016_/X VGND VGND VPWR VPWR _13017_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10229_ _09541_/B _09293_/B _08402_/X _10228_/Y VGND VGND VPWR VPWR _10230_/B sky130_fd_sc_hd__o22ai_2
X_14968_ _14984_/A _14984_/B _14967_/Y VGND VGND VPWR VPWR _14968_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14899_ _14812_/A _14812_/B _14812_/Y VGND VGND VPWR VPWR _14899_/X sky130_fd_sc_hd__a21o_1
X_13919_ _14627_/A _13846_/B _13846_/Y VGND VGND VPWR VPWR _13919_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09110_ _09717_/A _09113_/B VGND VGND VPWR VPWR _09110_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09041_ _09041_/A _09041_/B VGND VGND VPWR VPWR _09064_/A sky130_fd_sc_hd__or2_1
XFILLER_128_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09943_ _12932_/A VGND VGND VPWR VPWR _11843_/A sky130_fd_sc_hd__inv_2
XFILLER_58_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _08749_/Y _09873_/A _08749_/A _09937_/B VGND VGND VPWR VPWR _09874_/X sky130_fd_sc_hd__a22o_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _08825_/A VGND VGND VPWR VPWR _09252_/B sky130_fd_sc_hd__inv_2
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08756_ _09448_/A _09478_/B _08708_/Y VGND VGND VPWR VPWR _08757_/A sky130_fd_sc_hd__a21oi_2
XFILLER_26_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08687_ _09555_/A _08571_/A _08573_/Y _08686_/X VGND VGND VPWR VPWR _08687_/X sky130_fd_sc_hd__o22a_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09308_ _09286_/Y _09306_/Y _09307_/Y VGND VGND VPWR VPWR _09310_/B sky130_fd_sc_hd__o21ai_1
XFILLER_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10580_ _11867_/A _10651_/B _10579_/Y VGND VGND VPWR VPWR _10580_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09239_ _09539_/A _09687_/A _09230_/Y _09238_/Y VGND VGND VPWR VPWR _09239_/X sky130_fd_sc_hd__o22a_1
XFILLER_126_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12250_ _12249_/Y _12156_/X _12196_/Y VGND VGND VPWR VPWR _12250_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11201_ _13363_/A VGND VGND VPWR VPWR _14021_/A sky130_fd_sc_hd__inv_2
X_12181_ _12266_/B _12180_/X _12266_/B _12180_/X VGND VGND VPWR VPWR _12262_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11132_ _09993_/A _09993_/B _09993_/Y VGND VGND VPWR VPWR _11133_/A sky130_fd_sc_hd__o21ai_1
X_15940_ _15888_/A _15888_/B _15888_/Y VGND VGND VPWR VPWR _15940_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11063_ _13754_/A _11063_/B VGND VGND VPWR VPWR _13096_/A sky130_fd_sc_hd__or2_1
X_15871_ _15894_/A _15894_/B VGND VGND VPWR VPWR _15871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10014_ _10014_/A _10014_/B VGND VGND VPWR VPWR _10050_/B sky130_fd_sc_hd__nor2_1
X_14822_ _14794_/A _14794_/B _14794_/X _14821_/X VGND VGND VPWR VPWR _14822_/X sky130_fd_sc_hd__o22a_1
XFILLER_76_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11965_ _12038_/A _11963_/X _11964_/X VGND VGND VPWR VPWR _11965_/X sky130_fd_sc_hd__o21a_1
X_14753_ _12277_/Y _14752_/X _12277_/Y _14752_/X VGND VGND VPWR VPWR _14754_/B sky130_fd_sc_hd__o2bb2a_1
X_10916_ _14619_/A _10916_/B VGND VGND VPWR VPWR _10916_/X sky130_fd_sc_hd__or2_1
X_14684_ _14746_/A _14746_/B VGND VGND VPWR VPWR _14684_/Y sky130_fd_sc_hd__nand2_1
X_13704_ _13724_/A _13702_/X _13703_/X VGND VGND VPWR VPWR _13704_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16423_ _16468_/Q VGND VGND VPWR VPWR _16447_/A sky130_fd_sc_hd__inv_2
X_11896_ _11882_/Y _11894_/Y _11895_/Y VGND VGND VPWR VPWR _11897_/A sky130_fd_sc_hd__o21ai_2
X_13635_ _13593_/Y _13632_/Y _13634_/Y VGND VGND VPWR VPWR _13636_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10847_ _10847_/A VGND VGND VPWR VPWR _10847_/Y sky130_fd_sc_hd__inv_2
X_16354_ _16332_/A _16332_/B _16332_/Y VGND VGND VPWR VPWR _16354_/Y sky130_fd_sc_hd__o21ai_1
X_13566_ _15030_/A _13528_/B _13528_/Y VGND VGND VPWR VPWR _13566_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10778_ _09657_/X _10777_/X _09657_/X _10777_/X VGND VGND VPWR VPWR _10779_/B sky130_fd_sc_hd__a2bb2oi_1
X_16285_ _16268_/A _16334_/A _16268_/Y VGND VGND VPWR VPWR _16285_/Y sky130_fd_sc_hd__o21ai_1
X_12517_ _12517_/A _12517_/B VGND VGND VPWR VPWR _12517_/Y sky130_fd_sc_hd__nand2_1
X_15305_ _15345_/A _15345_/B VGND VGND VPWR VPWR _15369_/A sky130_fd_sc_hd__and2_1
X_13497_ _11536_/X _13492_/X _11536_/X _13492_/X VGND VGND VPWR VPWR _13498_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15236_ _15227_/X _15235_/Y _15227_/X _15235_/Y VGND VGND VPWR VPWR _15237_/B sky130_fd_sc_hd__a2bb2o_1
X_12448_ _13973_/A _12447_/B _12447_/Y VGND VGND VPWR VPWR _12448_/X sky130_fd_sc_hd__a21o_1
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15167_ _15167_/A _15167_/B VGND VGND VPWR VPWR _15167_/Y sky130_fd_sc_hd__nor2_1
X_12379_ _12379_/A _12379_/B VGND VGND VPWR VPWR _12379_/X sky130_fd_sc_hd__or2_1
XFILLER_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14118_ _14057_/X _14117_/X _14057_/X _14117_/X VGND VGND VPWR VPWR _14121_/A sky130_fd_sc_hd__a2bb2o_1
X_15098_ _15057_/A _15057_/B _15057_/Y _15097_/X VGND VGND VPWR VPWR _15098_/X sky130_fd_sc_hd__a2bb2o_1
X_14049_ _14815_/A _14048_/B _14047_/X _14048_/Y VGND VGND VPWR VPWR _14049_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08610_ _08610_/A _10113_/B VGND VGND VPWR VPWR _08611_/A sky130_fd_sc_hd__or2_1
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09590_ _09556_/X _09589_/X _09556_/X _09589_/X VGND VGND VPWR VPWR _09660_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08541_ _09529_/A VGND VGND VPWR VPWR _09472_/B sky130_fd_sc_hd__inv_2
XFILLER_63_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08472_ input3/X input19/X VGND VGND VPWR VPWR _08472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09024_ _08819_/A _08618_/X _09024_/S VGND VGND VPWR VPWR _09547_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09926_ _11298_/A _11297_/A VGND VGND VPWR VPWR _09926_/X sky130_fd_sc_hd__or2_1
XFILLER_131_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09857_ _09857_/A _09857_/B VGND VGND VPWR VPWR _09904_/A sky130_fd_sc_hd__or2_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08808_ _10127_/A VGND VGND VPWR VPWR _08810_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09788_ _09788_/A _09788_/B VGND VGND VPWR VPWR _09788_/X sky130_fd_sc_hd__or2_1
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08739_ _08739_/A VGND VGND VPWR VPWR _08739_/Y sky130_fd_sc_hd__inv_2
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11750_ _11750_/A _11750_/B VGND VGND VPWR VPWR _11750_/X sky130_fd_sc_hd__or2_1
XFILLER_121_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10701_ _11978_/A _10781_/B VGND VGND VPWR VPWR _10701_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11668_/A _15433_/A _11668_/Y _11573_/Y VGND VGND VPWR VPWR _11681_/Y sky130_fd_sc_hd__o2bb2ai_1
X_13420_ _13358_/X _13419_/X _13358_/X _13419_/X VGND VGND VPWR VPWR _13420_/Y sky130_fd_sc_hd__a2bb2oi_2
X_10632_ _10744_/A _10632_/B VGND VGND VPWR VPWR _10632_/Y sky130_fd_sc_hd__nand2_1
X_13351_ _13351_/A VGND VGND VPWR VPWR _15473_/A sky130_fd_sc_hd__buf_1
X_10563_ _10562_/A _10561_/Y _10562_/Y _10561_/A _10974_/A VGND VGND VPWR VPWR _10673_/B
+ sky130_fd_sc_hd__a221o_1
X_16070_ _16112_/A _16112_/B VGND VGND VPWR VPWR _16070_/X sky130_fd_sc_hd__and2_1
X_12302_ _12246_/X _12301_/Y _12246_/X _12301_/Y VGND VGND VPWR VPWR _12303_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13282_ _14729_/A _13282_/B VGND VGND VPWR VPWR _13282_/Y sky130_fd_sc_hd__nand2_1
X_10494_ _11839_/A VGND VGND VPWR VPWR _13621_/A sky130_fd_sc_hd__buf_1
X_15021_ _11751_/X _14999_/X _11751_/X _14999_/X VGND VGND VPWR VPWR _15032_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12233_ _12233_/A _12134_/X VGND VGND VPWR VPWR _12233_/X sky130_fd_sc_hd__or2b_1
XFILLER_107_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12164_ _12163_/Y _12072_/X _12095_/Y VGND VGND VPWR VPWR _12164_/X sky130_fd_sc_hd__o21a_1
X_11115_ _12160_/A _11115_/B VGND VGND VPWR VPWR _11115_/Y sky130_fd_sc_hd__nor2_1
X_12095_ _12095_/A _12163_/B VGND VGND VPWR VPWR _12095_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15923_ _15899_/X _15922_/Y _15899_/X _15922_/Y VGND VGND VPWR VPWR _15962_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11046_ _13922_/A _11081_/B VGND VGND VPWR VPWR _11228_/A sky130_fd_sc_hd__and2_1
XFILLER_77_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15854_ _12649_/Y _15853_/Y _14163_/B VGND VGND VPWR VPWR _15854_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15785_ _15785_/A _15667_/X VGND VGND VPWR VPWR _15785_/X sky130_fd_sc_hd__or2b_1
X_14805_ _14726_/Y _14804_/X _14726_/Y _14804_/X VGND VGND VPWR VPWR _14806_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14736_ _14788_/A _14734_/X _14735_/X VGND VGND VPWR VPWR _14736_/X sky130_fd_sc_hd__o21a_1
X_12997_ _13012_/A _13013_/B VGND VGND VPWR VPWR _13090_/A sky130_fd_sc_hd__and2_1
XFILLER_17_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11948_ _13078_/A _11970_/B VGND VGND VPWR VPWR _11948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14667_ _15240_/A VGND VGND VPWR VPWR _14746_/A sky130_fd_sc_hd__buf_1
X_11879_ _12990_/A _11898_/B VGND VGND VPWR VPWR _11879_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16406_ _16406_/A VGND VGND VPWR VPWR _16406_/Y sky130_fd_sc_hd__inv_2
X_13618_ _13610_/Y _13612_/Y _13617_/Y VGND VGND VPWR VPWR _13618_/X sky130_fd_sc_hd__o21a_1
X_14598_ _14597_/A _14597_/B _14597_/Y VGND VGND VPWR VPWR _14598_/X sky130_fd_sc_hd__a21o_1
X_16337_ _16284_/Y _16335_/X _16336_/Y VGND VGND VPWR VPWR _16337_/X sky130_fd_sc_hd__o21a_1
X_13549_ _13549_/A VGND VGND VPWR VPWR _13549_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16268_ _16268_/A _16268_/B VGND VGND VPWR VPWR _16268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16199_ _16104_/A _16104_/B _16104_/Y VGND VGND VPWR VPWR _16199_/X sky130_fd_sc_hd__o21a_1
XFILLER_114_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15219_ _15208_/A _15208_/B _15208_/Y _15218_/X VGND VGND VPWR VPWR _15219_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09711_ _09709_/A _09709_/B _09709_/Y _09954_/A VGND VGND VPWR VPWR _09713_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09642_ _09960_/A _09645_/B VGND VGND VPWR VPWR _09642_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09573_ _09559_/X _09572_/X _09559_/X _09572_/X VGND VGND VPWR VPWR _09666_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08524_/A VGND VGND VPWR VPWR _08524_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08455_ _08454_/A _08313_/Y _08454_/Y _08313_/A _08441_/X VGND VGND VPWR VPWR _08532_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08386_ _09228_/B VGND VGND VPWR VPWR _08386_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09007_ _08844_/A _09005_/Y _09006_/Y VGND VGND VPWR VPWR _09007_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09909_ _09734_/A _09904_/Y _09859_/B VGND VGND VPWR VPWR _09909_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12920_ _13003_/A _12920_/B VGND VGND VPWR VPWR _12920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12851_ _12807_/Y _12849_/X _12850_/Y VGND VGND VPWR VPWR _12851_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11802_ _11847_/A VGND VGND VPWR VPWR _12771_/A sky130_fd_sc_hd__buf_1
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15570_ _15655_/B VGND VGND VPWR VPWR _15571_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12732_/Y _12780_/X _12781_/Y VGND VGND VPWR VPWR _12782_/X sky130_fd_sc_hd__o21a_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14545_/A _14519_/X _14520_/X VGND VGND VPWR VPWR _14521_/X sky130_fd_sc_hd__o21a_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ _11733_/A _11733_/B VGND VGND VPWR VPWR _11733_/X sky130_fd_sc_hd__or2_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _13926_/A _14427_/B _13926_/A _14427_/B VGND VGND VPWR VPWR _14452_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11664_ _11664_/A _11664_/B VGND VGND VPWR VPWR _11664_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13403_ _13403_/A _13355_/X VGND VGND VPWR VPWR _13403_/X sky130_fd_sc_hd__or2b_1
X_10615_ _11889_/A VGND VGND VPWR VPWR _13001_/A sky130_fd_sc_hd__buf_1
XFILLER_128_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16122_ _16138_/A _16140_/A _16121_/X VGND VGND VPWR VPWR _16122_/X sky130_fd_sc_hd__o21a_1
X_14383_ _15636_/A _14381_/X _14382_/X VGND VGND VPWR VPWR _14383_/X sky130_fd_sc_hd__o21a_1
X_11595_ _11595_/A VGND VGND VPWR VPWR _11595_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13334_ _13334_/A _13334_/B VGND VGND VPWR VPWR _13334_/X sky130_fd_sc_hd__and2_1
XFILLER_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10546_ _09981_/A _09981_/B _09981_/Y VGND VGND VPWR VPWR _10547_/A sky130_fd_sc_hd__o21ai_1
X_16053_ _16053_/A _16053_/B VGND VGND VPWR VPWR _16062_/B sky130_fd_sc_hd__or2_1
XFILLER_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13265_ _14429_/A VGND VGND VPWR VPWR _13274_/A sky130_fd_sc_hd__clkbuf_2
X_10477_ _10452_/X _10476_/X _10452_/X _10476_/X VGND VGND VPWR VPWR _10544_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12216_ _12216_/A _12145_/X VGND VGND VPWR VPWR _12216_/X sky130_fd_sc_hd__or2b_1
X_15004_ _11926_/A _15003_/X _11925_/X VGND VGND VPWR VPWR _15004_/X sky130_fd_sc_hd__o21a_1
X_13196_ _13196_/A _13196_/B VGND VGND VPWR VPWR _13196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12147_ _13910_/A _12147_/B VGND VGND VPWR VPWR _12147_/X sky130_fd_sc_hd__or2_1
X_12078_ _12078_/A VGND VGND VPWR VPWR _12167_/A sky130_fd_sc_hd__inv_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15906_ _15906_/A _15906_/B VGND VGND VPWR VPWR _15906_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11029_ _13556_/A VGND VGND VPWR VPWR _12846_/A sky130_fd_sc_hd__buf_1
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15837_ _16136_/A VGND VGND VPWR VPWR _16277_/A sky130_fd_sc_hd__inv_2
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15768_ _15778_/B _15768_/B VGND VGND VPWR VPWR _15787_/A sky130_fd_sc_hd__or2_1
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15699_ _15553_/Y _15698_/X _15553_/Y _15698_/X VGND VGND VPWR VPWR _15700_/B sky130_fd_sc_hd__a2bb2oi_1
X_14719_ _14644_/A _14644_/B _14644_/Y VGND VGND VPWR VPWR _14719_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08240_ input6/X VGND VGND VPWR VPWR _08306_/B sky130_fd_sc_hd__inv_2
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09625_ _09503_/A _09505_/Y _09503_/Y VGND VGND VPWR VPWR _09625_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09556_ _09595_/A _09554_/X _09595_/B VGND VGND VPWR VPWR _09556_/X sky130_fd_sc_hd__o21ba_1
XFILLER_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09487_ _08781_/A _09471_/X _08781_/A _09471_/X VGND VGND VPWR VPWR _09488_/B sky130_fd_sc_hd__o2bb2a_1
X_08507_ _08662_/A _09677_/B VGND VGND VPWR VPWR _08509_/A sky130_fd_sc_hd__or2_4
XFILLER_51_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08438_ _08565_/B _08433_/X _09452_/A VGND VGND VPWR VPWR _08439_/A sky130_fd_sc_hd__o21ai_1
X_08369_ _08266_/A input13/X _08347_/B _08414_/A VGND VGND VPWR VPWR _08418_/A sky130_fd_sc_hd__o22a_1
X_11380_ _11391_/A _11380_/B VGND VGND VPWR VPWR _12312_/A sky130_fd_sc_hd__or2_1
X_10400_ _11775_/A _10400_/B VGND VGND VPWR VPWR _10400_/X sky130_fd_sc_hd__and2_1
XFILLER_109_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10331_ _09954_/A _10330_/A _09954_/Y _10330_/Y _10446_/A VGND VGND VPWR VPWR _11719_/A
+ sky130_fd_sc_hd__o221a_1
X_13050_ _13050_/A _13030_/X VGND VGND VPWR VPWR _13050_/X sky130_fd_sc_hd__or2b_1
XFILLER_3_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10262_ _09377_/B _10239_/B _10239_/X _11329_/A VGND VGND VPWR VPWR _11533_/A sky130_fd_sc_hd__a22o_1
X_12001_ _12777_/A _12076_/A _12000_/Y VGND VGND VPWR VPWR _12001_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10193_ _10194_/A _10194_/B VGND VGND VPWR VPWR _10193_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13952_ _15410_/A _13952_/B VGND VGND VPWR VPWR _13952_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12903_ _14463_/A _12928_/B VGND VGND VPWR VPWR _12903_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13883_ _13883_/A _13883_/B VGND VGND VPWR VPWR _13883_/X sky130_fd_sc_hd__or2_1
XFILLER_62_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15622_ _15675_/A _15675_/B VGND VGND VPWR VPWR _15622_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12834_ _10422_/A _12830_/X _10426_/A _12833_/Y VGND VGND VPWR VPWR _12836_/B sky130_fd_sc_hd__o22a_1
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15491_/X _15551_/X _15573_/B VGND VGND VPWR VPWR _15553_/Y sky130_fd_sc_hd__o21ai_2
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12765_ _12765_/A _12765_/B VGND VGND VPWR VPWR _12765_/Y sky130_fd_sc_hd__nand2_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _15211_/A _14510_/B VGND VGND VPWR VPWR _14565_/A sky130_fd_sc_hd__and2_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11716_/A VGND VGND VPWR VPWR _11717_/B sky130_fd_sc_hd__inv_2
X_15484_ _14778_/A _15443_/B _15443_/X _15483_/X VGND VGND VPWR VPWR _15484_/X sky130_fd_sc_hd__o22a_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A _12696_/B VGND VGND VPWR VPWR _12696_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11647_ _12443_/A _11647_/B VGND VGND VPWR VPWR _11647_/X sky130_fd_sc_hd__or2_1
X_14435_ _14423_/A _14423_/B _14423_/Y _14434_/X VGND VGND VPWR VPWR _14435_/X sky130_fd_sc_hd__o2bb2a_1
Xinput13 wbs_adr_i[5] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_1
XFILLER_30_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput24 wbs_dat_i[15] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_2
XFILLER_128_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14366_ _14366_/A VGND VGND VPWR VPWR _14366_/Y sky130_fd_sc_hd__inv_2
X_11578_ _11629_/A VGND VGND VPWR VPWR _13133_/A sky130_fd_sc_hd__buf_1
X_16105_ _16101_/Y _16103_/X _16104_/Y VGND VGND VPWR VPWR _16105_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13317_ _14741_/A _13300_/B _13300_/Y VGND VGND VPWR VPWR _13317_/Y sky130_fd_sc_hd__o21ai_1
X_10529_ _11839_/A _10529_/B VGND VGND VPWR VPWR _10529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16036_ _16036_/A _16036_/B VGND VGND VPWR VPWR _16036_/Y sky130_fd_sc_hd__nand2_1
X_14297_ _15972_/A _14403_/B VGND VGND VPWR VPWR _14297_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13248_ _13192_/A _13192_/B _13192_/Y VGND VGND VPWR VPWR _13248_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_97_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13179_ _13833_/A VGND VGND VPWR VPWR _15329_/A sky130_fd_sc_hd__buf_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09410_ _09409_/A _09409_/B _10402_/A _09409_/Y VGND VGND VPWR VPWR _09412_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_53_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09341_ _09341_/A _09341_/B VGND VGND VPWR VPWR _09342_/B sky130_fd_sc_hd__or2_1
XFILLER_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09272_ _09272_/A VGND VGND VPWR VPWR _09275_/A sky130_fd_sc_hd__inv_2
XFILLER_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08987_ _08870_/Y _08985_/X _08986_/Y VGND VGND VPWR VPWR _08987_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10880_ _10883_/A VGND VGND VPWR VPWR _14631_/A sky130_fd_sc_hd__buf_1
XFILLER_73_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09608_ _09550_/X _09607_/Y _09550_/X _09607_/Y VGND VGND VPWR VPWR _09654_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09539_ _09539_/A _09539_/B VGND VGND VPWR VPWR _09539_/X sky130_fd_sc_hd__or2_1
XFILLER_71_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12550_ _14916_/A _12349_/B _12349_/Y VGND VGND VPWR VPWR _12551_/A sky130_fd_sc_hd__o21ai_1
X_12481_ _15556_/A _12452_/B _12452_/Y _12480_/Y VGND VGND VPWR VPWR _12481_/X sky130_fd_sc_hd__o2bb2a_1
X_11501_ _09929_/Y _11500_/X _09931_/A _09930_/Y _10792_/X VGND VGND VPWR VPWR _12946_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14220_ _14220_/A _12621_/X VGND VGND VPWR VPWR _14220_/X sky130_fd_sc_hd__or2b_1
X_11432_ _12224_/A _11230_/B _11230_/Y VGND VGND VPWR VPWR _11432_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14151_ _13969_/A _13970_/Y _13968_/X VGND VGND VPWR VPWR _14151_/X sky130_fd_sc_hd__o21a_1
XFILLER_125_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11363_ _12303_/A _11363_/B VGND VGND VPWR VPWR _11363_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13102_ _13096_/X _13100_/Y _13101_/Y VGND VGND VPWR VPWR _13102_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14082_ _14082_/A _14082_/B VGND VGND VPWR VPWR _14082_/Y sky130_fd_sc_hd__nor2_1
X_11294_ _12362_/A VGND VGND VPWR VPWR _13793_/A sky130_fd_sc_hd__buf_1
X_10314_ _10248_/A _10313_/A _10248_/Y _10313_/Y _10472_/A VGND VGND VPWR VPWR _11757_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13033_ _13045_/A _13031_/X _13032_/X VGND VGND VPWR VPWR _13033_/X sky130_fd_sc_hd__o21a_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ _10245_/A VGND VGND VPWR VPWR _10247_/A sky130_fd_sc_hd__inv_2
XFILLER_121_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10176_ _10123_/A _10123_/B _10124_/B VGND VGND VPWR VPWR _10180_/A sky130_fd_sc_hd__a21bo_1
XFILLER_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14984_ _14984_/A _14984_/B VGND VGND VPWR VPWR _14984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13935_ _10906_/A _13934_/Y _10906_/A _13934_/Y VGND VGND VPWR VPWR _13938_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13866_ _13864_/Y _13865_/Y _13789_/Y VGND VGND VPWR VPWR _13866_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15605_ _15605_/A _14390_/X VGND VGND VPWR VPWR _15605_/X sky130_fd_sc_hd__or2b_1
XFILLER_74_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12817_ _12767_/A _12767_/B _12767_/Y VGND VGND VPWR VPWR _12817_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13797_ _13797_/A _13797_/B VGND VGND VPWR VPWR _13797_/X sky130_fd_sc_hd__or2_1
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15536_ _15540_/A _15540_/B VGND VGND VPWR VPWR _15536_/Y sky130_fd_sc_hd__nor2_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12748_ _12698_/A _12698_/B _12698_/Y VGND VGND VPWR VPWR _12748_/X sky130_fd_sc_hd__a21o_1
X_15467_ _15467_/A _15467_/B VGND VGND VPWR VPWR _15467_/Y sky130_fd_sc_hd__nand2_1
X_12679_ _12679_/A _12679_/B VGND VGND VPWR VPWR _12679_/Y sky130_fd_sc_hd__nor2_1
X_14418_ _15032_/A _11753_/Y _11772_/Y _14417_/X VGND VGND VPWR VPWR _14418_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15398_ _15398_/A _15398_/B VGND VGND VPWR VPWR _15398_/X sky130_fd_sc_hd__or2_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14349_ _15878_/A _14254_/B _14254_/Y VGND VGND VPWR VPWR _14349_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16019_ _16034_/A _16034_/B VGND VGND VPWR VPWR _16019_/Y sky130_fd_sc_hd__nor2_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _09888_/A _09888_/B _09888_/X VGND VGND VPWR VPWR _09928_/A sky130_fd_sc_hd__a21bo_1
X_08910_ _08819_/A _10126_/A _08819_/Y VGND VGND VPWR VPWR _08910_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08944_/B VGND VGND VPWR VPWR _10123_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _09332_/A _09474_/B _08710_/Y VGND VGND VPWR VPWR _08773_/A sky130_fd_sc_hd__a21oi_2
XFILLER_38_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09324_ _09324_/A _10129_/A VGND VGND VPWR VPWR _10047_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09255_ _09459_/A _10123_/A _08944_/X _09301_/A VGND VGND VPWR VPWR _09255_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_21_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09186_ _09182_/Y _09184_/Y _09185_/Y VGND VGND VPWR VPWR _09191_/B sky130_fd_sc_hd__o21ai_1
XFILLER_119_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10030_ _10035_/B _10029_/X _10035_/A VGND VGND VPWR VPWR _10030_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_102_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11981_ _13637_/A _11981_/B VGND VGND VPWR VPWR _11981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13720_ _13720_/A _13720_/B VGND VGND VPWR VPWR _13720_/X sky130_fd_sc_hd__or2_1
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10932_ _09659_/X _10931_/X _09659_/X _10931_/X VGND VGND VPWR VPWR _10933_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_29_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10863_ _12057_/A VGND VGND VPWR VPWR _10867_/A sky130_fd_sc_hd__inv_2
X_13651_ _13646_/X _13650_/Y _13646_/X _13650_/Y VGND VGND VPWR VPWR _13706_/B sky130_fd_sc_hd__a2bb2o_1
X_16370_ _16323_/X _16369_/Y _16323_/X _16369_/Y VGND VGND VPWR VPWR _16397_/D sky130_fd_sc_hd__a2bb2o_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12602_ _12602_/A VGND VGND VPWR VPWR _12602_/Y sky130_fd_sc_hd__inv_2
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10794_ _12938_/A VGND VGND VPWR VPWR _12005_/A sky130_fd_sc_hd__inv_2
X_13582_ _15042_/A _13510_/B _13510_/Y VGND VGND VPWR VPWR _13582_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ _12533_/A _12533_/B VGND VGND VPWR VPWR _12533_/Y sky130_fd_sc_hd__nand2_1
X_15321_ _14576_/A _15264_/B _15264_/Y VGND VGND VPWR VPWR _15321_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15252_ _15252_/A _15252_/B VGND VGND VPWR VPWR _15252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14203_ _12626_/X _14202_/X _12626_/X _14202_/X VGND VGND VPWR VPWR _14266_/B sky130_fd_sc_hd__a2bb2o_1
X_12464_ _13989_/A _12466_/B VGND VGND VPWR VPWR _12474_/A sky130_fd_sc_hd__and2_1
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11415_ _14047_/A _13350_/A VGND VGND VPWR VPWR _13406_/B sky130_fd_sc_hd__or2_1
X_12395_ _12361_/Y _12394_/X _12361_/Y _12394_/X VGND VGND VPWR VPWR _12397_/B sky130_fd_sc_hd__o2bb2a_1
X_15183_ _15156_/X _15182_/Y _15156_/X _15182_/Y VGND VGND VPWR VPWR _15184_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14134_ _14128_/X _14131_/Y _14868_/A _14133_/Y VGND VGND VPWR VPWR _14134_/X sky130_fd_sc_hd__o22a_1
X_11346_ _11283_/X _11345_/Y _11283_/X _11345_/Y VGND VGND VPWR VPWR _11480_/B sky130_fd_sc_hd__o2bb2a_1
X_14065_ _14135_/A _14063_/X _14064_/X VGND VGND VPWR VPWR _14065_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11277_ _11276_/A _11276_/B _11276_/X _11103_/X VGND VGND VPWR VPWR _11277_/X sky130_fd_sc_hd__o22a_1
X_13016_ _14493_/A _13016_/B VGND VGND VPWR VPWR _13016_/X sky130_fd_sc_hd__or2_1
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10228_ _10228_/A _10228_/B VGND VGND VPWR VPWR _10228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10159_ _10159_/A _10159_/B VGND VGND VPWR VPWR _10159_/Y sky130_fd_sc_hd__nor2_1
X_14967_ _14984_/A _14984_/B VGND VGND VPWR VPWR _14967_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14898_ _14908_/A _14908_/B VGND VGND VPWR VPWR _14898_/Y sky130_fd_sc_hd__nor2_1
X_13918_ _13918_/A VGND VGND VPWR VPWR _15404_/A sky130_fd_sc_hd__buf_1
XFILLER_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13849_ _13818_/Y _13847_/X _13848_/Y VGND VGND VPWR VPWR _13849_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15519_ _15519_/A _15519_/B VGND VGND VPWR VPWR _15519_/X sky130_fd_sc_hd__or2_1
X_09040_ _09040_/A VGND VGND VPWR VPWR _09040_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09942_ _09806_/Y _09854_/Y _09897_/A _09855_/X _10792_/A VGND VGND VPWR VPWR _12932_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09873_ _09873_/A VGND VGND VPWR VPWR _09937_/B sky130_fd_sc_hd__inv_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08823_/X _08726_/X _08823_/A _08726_/X VGND VGND VPWR VPWR _08825_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08755_ _08755_/A VGND VGND VPWR VPWR _09478_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08686_ _09553_/A _08584_/A _08586_/Y _08685_/X VGND VGND VPWR VPWR _08686_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09307_ _10245_/A _09307_/B VGND VGND VPWR VPWR _09307_/Y sky130_fd_sc_hd__nand2_1
X_09238_ _09238_/A VGND VGND VPWR VPWR _09238_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09169_ _09169_/A VGND VGND VPWR VPWR _09750_/A sky130_fd_sc_hd__inv_2
X_12180_ _12180_/A _12179_/X VGND VGND VPWR VPWR _12180_/X sky130_fd_sc_hd__or2b_1
X_11200_ _09130_/Y _11199_/A _09130_/A _11199_/Y _11219_/B VGND VGND VPWR VPWR _13363_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11131_ _13507_/A _11130_/B _11130_/X _10954_/X VGND VGND VPWR VPWR _11131_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11062_ _11062_/A VGND VGND VPWR VPWR _11064_/B sky130_fd_sc_hd__buf_1
X_15870_ _14208_/X _15844_/X _14208_/X _15844_/X VGND VGND VPWR VPWR _15894_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10013_ _10013_/A _10013_/B VGND VGND VPWR VPWR _10047_/B sky130_fd_sc_hd__nor2_1
X_14821_ _14798_/A _14798_/B _14798_/X _14820_/X VGND VGND VPWR VPWR _14821_/X sky130_fd_sc_hd__o22a_1
XFILLER_95_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11964_ _11964_/A _11964_/B VGND VGND VPWR VPWR _11964_/X sky130_fd_sc_hd__or2_1
XFILLER_56_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14752_ _15046_/A _12262_/Y _12182_/Y _14672_/X VGND VGND VPWR VPWR _14752_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10915_ _10915_/A VGND VGND VPWR VPWR _14619_/A sky130_fd_sc_hd__buf_1
X_14683_ _14668_/X _14682_/X _14668_/X _14682_/X VGND VGND VPWR VPWR _14746_/B sky130_fd_sc_hd__a2bb2o_1
X_11895_ _12994_/A _11895_/B VGND VGND VPWR VPWR _11895_/Y sky130_fd_sc_hd__nand2_1
X_13703_ _13703_/A _13703_/B VGND VGND VPWR VPWR _13703_/X sky130_fd_sc_hd__or2_1
XFILLER_32_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16422_ _16474_/Q _16473_/Q VGND VGND VPWR VPWR _16447_/B sky130_fd_sc_hd__or2_1
X_13634_ _15128_/A _13634_/B VGND VGND VPWR VPWR _13634_/Y sky130_fd_sc_hd__nand2_1
X_10846_ _09424_/A _09424_/B _09424_/Y VGND VGND VPWR VPWR _10847_/A sky130_fd_sc_hd__o21ai_1
X_16353_ _08230_/X _16467_/Q _08233_/X _16402_/A _16343_/X VGND VGND VPWR VPWR _16467_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15304_ _15279_/X _15303_/Y _15279_/X _15303_/Y VGND VGND VPWR VPWR _15345_/B sky130_fd_sc_hd__a2bb2o_1
X_13565_ _13565_/A VGND VGND VPWR VPWR _13565_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10777_ _09987_/A _09658_/B _09658_/Y VGND VGND VPWR VPWR _10777_/X sky130_fd_sc_hd__o21a_1
X_16284_ _16336_/A _16336_/B VGND VGND VPWR VPWR _16284_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12516_ _13444_/A _12303_/B _12303_/Y VGND VGND VPWR VPWR _12517_/B sky130_fd_sc_hd__o21a_1
X_13496_ _13496_/A VGND VGND VPWR VPWR _15104_/A sky130_fd_sc_hd__buf_1
XFILLER_117_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15235_ _15181_/A _15181_/B _15181_/Y VGND VGND VPWR VPWR _15235_/Y sky130_fd_sc_hd__o21ai_1
X_12447_ _13973_/A _12447_/B VGND VGND VPWR VPWR _12447_/Y sky130_fd_sc_hd__nor2_1
X_15166_ _15164_/X _15165_/Y _15164_/X _15165_/Y VGND VGND VPWR VPWR _15167_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14117_ _14117_/A _14058_/X VGND VGND VPWR VPWR _14117_/X sky130_fd_sc_hd__or2b_1
X_12378_ _12379_/A _12379_/B VGND VGND VPWR VPWR _12380_/A sky130_fd_sc_hd__and2_1
XFILLER_125_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15097_ _15060_/A _15060_/B _15060_/Y _15096_/X VGND VGND VPWR VPWR _15097_/X sky130_fd_sc_hd__a2bb2o_1
X_11329_ _11329_/A _11329_/B VGND VGND VPWR VPWR _11329_/Y sky130_fd_sc_hd__nand2_1
X_14048_ _14048_/A _14048_/B VGND VGND VPWR VPWR _14048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15999_ _15999_/A _15964_/X VGND VGND VPWR VPWR _15999_/X sky130_fd_sc_hd__or2b_1
XFILLER_94_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08540_ _08701_/A _08540_/B VGND VGND VPWR VPWR _09529_/A sky130_fd_sc_hd__or2_2
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08471_ input4/X input20/X VGND VGND VPWR VPWR _08471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09023_ _08605_/X _08904_/X _09023_/S VGND VGND VPWR VPWR _09549_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09925_ _09861_/A _09861_/B _09924_/Y VGND VGND VPWR VPWR _11297_/A sky130_fd_sc_hd__a21oi_1
XFILLER_112_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09856_ _09856_/A _09856_/B VGND VGND VPWR VPWR _09857_/B sky130_fd_sc_hd__or2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08807_ _08806_/A _08729_/A _08806_/Y _08729_/Y VGND VGND VPWR VPWR _10127_/A sky130_fd_sc_hd__o22a_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09787_ _09788_/A _09788_/B VGND VGND VPWR VPWR _11494_/A sky130_fd_sc_hd__and2_1
X_08738_ _08711_/Y _08736_/Y _08737_/X VGND VGND VPWR VPWR _08739_/A sky130_fd_sc_hd__o21ai_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08669_ _09541_/B VGND VGND VPWR VPWR _10228_/A sky130_fd_sc_hd__inv_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10652_/X _10699_/Y _10652_/X _10699_/Y VGND VGND VPWR VPWR _10781_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11678_/Y _11679_/X _11678_/Y _11679_/X VGND VGND VPWR VPWR _11680_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10631_ _10631_/A VGND VGND VPWR VPWR _10631_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13350_ _13350_/A VGND VGND VPWR VPWR _13350_/Y sky130_fd_sc_hd__inv_2
X_10562_ _10562_/A VGND VGND VPWR VPWR _10562_/Y sky130_fd_sc_hd__inv_2
X_12301_ _14012_/A _12203_/B _12203_/Y VGND VGND VPWR VPWR _12301_/Y sky130_fd_sc_hd__o21ai_1
X_13281_ _13281_/A VGND VGND VPWR VPWR _13281_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12232_ _12232_/A _12232_/B VGND VGND VPWR VPWR _12232_/Y sky130_fd_sc_hd__nor2_1
X_10493_ _12928_/A VGND VGND VPWR VPWR _11839_/A sky130_fd_sc_hd__inv_2
X_15020_ _15034_/A _15034_/B VGND VGND VPWR VPWR _15073_/A sky130_fd_sc_hd__and2_1
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12163_ _13706_/A _12163_/B VGND VGND VPWR VPWR _12163_/Y sky130_fd_sc_hd__nor2_1
X_11114_ _12252_/A VGND VGND VPWR VPWR _13048_/A sky130_fd_sc_hd__buf_1
X_12094_ _12074_/X _12093_/X _12074_/X _12093_/X VGND VGND VPWR VPWR _12163_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15922_ _15900_/A _15900_/B _15900_/Y VGND VGND VPWR VPWR _15922_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11045_ _10911_/X _11044_/X _10911_/X _11044_/X VGND VGND VPWR VPWR _11081_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15853_ _15853_/A VGND VGND VPWR VPWR _15853_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15784_ _15787_/A _15788_/B VGND VGND VPWR VPWR _15784_/Y sky130_fd_sc_hd__nor2_1
X_14804_ _14804_/A _14727_/X VGND VGND VPWR VPWR _14804_/X sky130_fd_sc_hd__or2b_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12996_ _12925_/X _12995_/Y _12925_/X _12995_/Y VGND VGND VPWR VPWR _13013_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14735_ _14735_/A _14735_/B VGND VGND VPWR VPWR _14735_/X sky130_fd_sc_hd__or2_1
X_11947_ _11900_/A _11946_/Y _11900_/A _11946_/Y VGND VGND VPWR VPWR _11970_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14666_ _14589_/X _14665_/Y _14607_/Y VGND VGND VPWR VPWR _14666_/X sky130_fd_sc_hd__o21a_1
X_11878_ _11838_/X _11877_/Y _11838_/X _11877_/Y VGND VGND VPWR VPWR _11898_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16405_ _16399_/Y _16400_/Y _16394_/Y _16393_/Y VGND VGND VPWR VPWR _16406_/A sky130_fd_sc_hd__a31o_1
X_13617_ _13003_/A _13616_/Y _12919_/A VGND VGND VPWR VPWR _13617_/Y sky130_fd_sc_hd__o21ai_1
X_14597_ _14597_/A _14597_/B VGND VGND VPWR VPWR _14597_/Y sky130_fd_sc_hd__nor2_1
X_10829_ _10962_/A _12080_/A VGND VGND VPWR VPWR _10829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16336_ _16336_/A _16336_/B VGND VGND VPWR VPWR _16336_/Y sky130_fd_sc_hd__nand2_1
X_13548_ _13548_/A _13548_/B VGND VGND VPWR VPWR _13549_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16267_ _16170_/Y _16265_/X _16266_/Y VGND VGND VPWR VPWR _16267_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15218_ _15211_/A _15211_/B _15211_/Y _15217_/X VGND VGND VPWR VPWR _15218_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13479_ _13479_/A _13479_/B VGND VGND VPWR VPWR _13479_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16198_ _16197_/A _16196_/Y _16197_/Y _16196_/A _15832_/A VGND VGND VPWR VPWR _16257_/A
+ sky130_fd_sc_hd__a221o_1
X_15149_ _15140_/A _15140_/B _15140_/Y _15148_/X VGND VGND VPWR VPWR _15149_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09710_ _09683_/A _09683_/B _09686_/A VGND VGND VPWR VPWR _09954_/A sky130_fd_sc_hd__a21bo_1
XFILLER_68_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09641_ _09637_/Y _10740_/A _09640_/Y VGND VGND VPWR VPWR _09645_/B sky130_fd_sc_hd__o21ai_1
X_09572_ _08694_/A _09152_/A _09526_/A VGND VGND VPWR VPWR _09572_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08523_ _09348_/B _09791_/C VGND VGND VPWR VPWR _08524_/A sky130_fd_sc_hd__or2_1
XFILLER_35_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08454_ _08454_/A VGND VGND VPWR VPWR _08454_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08385_ _08365_/Y _08384_/A _08365_/A _08384_/Y _08303_/A VGND VGND VPWR VPWR _09228_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09006_ _09006_/A VGND VGND VPWR VPWR _09006_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09908_ _09908_/A _09908_/B VGND VGND VPWR VPWR _09911_/A sky130_fd_sc_hd__and2_1
XFILLER_58_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09839_ _09839_/A VGND VGND VPWR VPWR _09839_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12850_ _12850_/A _12850_/B VGND VGND VPWR VPWR _12850_/Y sky130_fd_sc_hd__nand2_1
X_11801_ _11801_/A VGND VGND VPWR VPWR _11847_/A sky130_fd_sc_hd__inv_2
XFILLER_27_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _15196_/A _14520_/B VGND VGND VPWR VPWR _14520_/X sky130_fd_sc_hd__or2_1
X_12781_ _12781_/A _12781_/B VGND VGND VPWR VPWR _12781_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11731_/A _11731_/B _11730_/Y _11731_/Y VGND VGND VPWR VPWR _11742_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14463_/A _14463_/B VGND VGND VPWR VPWR _14451_/Y sky130_fd_sc_hd__nor2_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _11663_/A VGND VGND VPWR VPWR _11663_/Y sky130_fd_sc_hd__inv_2
X_14382_ _14382_/A _15952_/A VGND VGND VPWR VPWR _14382_/X sky130_fd_sc_hd__or2_1
X_13402_ _13405_/A VGND VGND VPWR VPWR _14904_/A sky130_fd_sc_hd__buf_1
X_10614_ _10618_/A _10756_/B VGND VGND VPWR VPWR _11889_/A sky130_fd_sc_hd__or2b_1
XFILLER_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16121_ _16121_/A _16121_/B VGND VGND VPWR VPWR _16121_/X sky130_fd_sc_hd__or2_1
X_13333_ _13284_/A _13332_/Y _13284_/A _13332_/Y VGND VGND VPWR VPWR _13334_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11594_ _09569_/A _09999_/B _10000_/A VGND VGND VPWR VPWR _11595_/A sky130_fd_sc_hd__o21ai_1
XFILLER_10_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10545_ _13519_/A _10544_/B _10544_/X _10443_/X VGND VGND VPWR VPWR _10545_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16052_ _16048_/Y _16050_/X _16051_/Y VGND VGND VPWR VPWR _16052_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13264_ _14725_/A _13276_/B VGND VGND VPWR VPWR _13264_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10476_ _10552_/A _12696_/A _10475_/Y VGND VGND VPWR VPWR _10476_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12215_ _12215_/A _12215_/B VGND VGND VPWR VPWR _12215_/Y sky130_fd_sc_hd__nand2_1
X_13195_ _13162_/Y _13193_/X _13194_/Y VGND VGND VPWR VPWR _13195_/X sky130_fd_sc_hd__o21a_1
X_15003_ _11860_/A _15002_/X _11859_/X VGND VGND VPWR VPWR _15003_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12146_ _12216_/A _12144_/X _12145_/X VGND VGND VPWR VPWR _12146_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12077_ _12075_/A _12075_/B _12075_/X _12076_/Y VGND VGND VPWR VPWR _12167_/B sky130_fd_sc_hd__a22o_1
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15905_ _14178_/X _15849_/X _14178_/X _15849_/X VGND VGND VPWR VPWR _15905_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11028_ _11028_/A VGND VGND VPWR VPWR _13556_/A sky130_fd_sc_hd__buf_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15836_ _16160_/A _15836_/B VGND VGND VPWR VPWR _16136_/A sky130_fd_sc_hd__or2_1
XFILLER_77_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15767_ _14905_/X _15766_/X _14905_/X _15766_/X VGND VGND VPWR VPWR _15768_/B sky130_fd_sc_hd__a2bb2oi_1
X_12979_ _14469_/A _12934_/B _12934_/Y VGND VGND VPWR VPWR _12979_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15698_ _14984_/A _15554_/B _15554_/Y VGND VGND VPWR VPWR _15698_/X sky130_fd_sc_hd__o21a_1
X_14718_ _15398_/A _14718_/B VGND VGND VPWR VPWR _14718_/X sky130_fd_sc_hd__and2_1
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14649_ _14638_/Y _14647_/Y _14648_/Y VGND VGND VPWR VPWR _14649_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16319_ _16311_/Y _16317_/X _16318_/Y VGND VGND VPWR VPWR _16319_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09624_ _09957_/A VGND VGND VPWR VPWR _09958_/A sky130_fd_sc_hd__buf_1
XFILLER_71_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09555_ _09555_/A _09555_/B VGND VGND VPWR VPWR _09595_/B sky130_fd_sc_hd__and2_1
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08506_ _08508_/A VGND VGND VPWR VPWR _09863_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09486_ _09486_/A _09486_/B VGND VGND VPWR VPWR _09486_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08437_ _08712_/A VGND VGND VPWR VPWR _09452_/A sky130_fd_sc_hd__buf_1
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08368_ _08269_/A input12/X _08353_/B _08409_/A VGND VGND VPWR VPWR _08414_/A sky130_fd_sc_hd__o22a_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08299_ _08237_/A input23/X _08238_/A _08296_/A VGND VGND VPWR VPWR _08299_/X sky130_fd_sc_hd__o22a_2
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10330_ _10330_/A VGND VGND VPWR VPWR _10330_/Y sky130_fd_sc_hd__inv_2
X_10261_ _09383_/B _10240_/B _10240_/X _11155_/A VGND VGND VPWR VPWR _11329_/A sky130_fd_sc_hd__a22o_1
XFILLER_105_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12000_ _12777_/A _12076_/A VGND VGND VPWR VPWR _12000_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10192_ _10238_/B _10139_/B _10139_/Y _10191_/X VGND VGND VPWR VPWR _10194_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_120_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13951_ _13913_/Y _13949_/X _13950_/Y VGND VGND VPWR VPWR _13951_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12902_ _12841_/X _12901_/Y _12841_/X _12901_/Y VGND VGND VPWR VPWR _12928_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13882_ _13883_/A _13883_/B VGND VGND VPWR VPWR _13884_/A sky130_fd_sc_hd__and2_1
XFILLER_19_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _14385_/X _15620_/X _14385_/X _15620_/X VGND VGND VPWR VPWR _15675_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12833_ _12832_/A _12832_/B _12832_/Y VGND VGND VPWR VPWR _12833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15552_/A _15552_/B VGND VGND VPWR VPWR _15573_/B sky130_fd_sc_hd__or2_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12760_/Y _12762_/Y _12763_/Y VGND VGND VPWR VPWR _12764_/X sky130_fd_sc_hd__o21a_1
X_15483_ _14782_/A _15446_/B _15446_/X _15482_/X VGND VGND VPWR VPWR _15483_/X sky130_fd_sc_hd__o22a_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _14458_/Y _14502_/X _14458_/Y _14502_/X VGND VGND VPWR VPWR _14510_/B sky130_fd_sc_hd__o2bb2a_1
X_11715_ _11715_/A VGND VGND VPWR VPWR _11788_/A sky130_fd_sc_hd__inv_2
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12695_ _10467_/A _12662_/A _10467_/Y _12662_/Y VGND VGND VPWR VPWR _12696_/B sky130_fd_sc_hd__o22a_1
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11646_ _12443_/A _11647_/B VGND VGND VPWR VPWR _11648_/A sky130_fd_sc_hd__and2_1
X_14434_ _14425_/A _14425_/B _14425_/Y _14433_/X VGND VGND VPWR VPWR _14434_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput14 wbs_adr_i[6] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_4
X_14365_ _14904_/A _13405_/B _13405_/X VGND VGND VPWR VPWR _14366_/A sky130_fd_sc_hd__o21ba_1
Xinput25 wbs_dat_i[1] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_4
X_11577_ _11576_/A _11576_/B _11576_/Y _09393_/X VGND VGND VPWR VPWR _11629_/A sky130_fd_sc_hd__o211a_1
XFILLER_128_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16104_ _16104_/A _16104_/B VGND VGND VPWR VPWR _16104_/Y sky130_fd_sc_hd__nand2_1
X_14296_ _14287_/X _14295_/X _14287_/X _14295_/X VGND VGND VPWR VPWR _14403_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13316_ _13371_/A _13371_/B VGND VGND VPWR VPWR _13379_/A sky130_fd_sc_hd__and2_1
X_10528_ _10506_/Y _10526_/X _10527_/Y VGND VGND VPWR VPWR _10528_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16035_ _16019_/Y _16033_/X _16034_/Y VGND VGND VPWR VPWR _16035_/X sky130_fd_sc_hd__o21a_1
X_13247_ _14421_/A VGND VGND VPWR VPWR _14731_/A sky130_fd_sc_hd__buf_1
X_10459_ _10459_/A VGND VGND VPWR VPWR _11854_/A sky130_fd_sc_hd__inv_2
XFILLER_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13178_ _15331_/A _13184_/B VGND VGND VPWR VPWR _13178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12129_ _12049_/A _12049_/B _12049_/Y VGND VGND VPWR VPWR _12129_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15819_ _16121_/A _15819_/B VGND VGND VPWR VPWR _16150_/B sky130_fd_sc_hd__or2_1
XFILLER_92_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09340_ _08753_/Y _09338_/Y _09339_/X VGND VGND VPWR VPWR _09340_/X sky130_fd_sc_hd__o21a_1
X_09271_ _09242_/X _09270_/X _09242_/X _09270_/X VGND VGND VPWR VPWR _09272_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08986_ _08986_/A _08986_/B VGND VGND VPWR VPWR _08986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09607_ _09607_/A _09607_/B VGND VGND VPWR VPWR _09607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09538_ _09538_/A _09538_/B VGND VGND VPWR VPWR _09538_/X sky130_fd_sc_hd__and2_1
X_11500_ _09928_/A _09928_/B _09931_/A VGND VGND VPWR VPWR _11500_/X sky130_fd_sc_hd__o21ba_1
X_09469_ _10013_/A _08572_/A _09453_/Y _09468_/X VGND VGND VPWR VPWR _09469_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12480_ _12480_/A VGND VGND VPWR VPWR _12480_/Y sky130_fd_sc_hd__inv_2
X_11431_ _12575_/A _11434_/B VGND VGND VPWR VPWR _11431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14150_ _14146_/X _14149_/Y _13450_/A _14149_/B VGND VGND VPWR VPWR _14150_/X sky130_fd_sc_hd__a2bb2o_1
X_11362_ _11260_/X _11361_/Y _11260_/X _11361_/Y VGND VGND VPWR VPWR _11363_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13101_ _13101_/A _13101_/B VGND VGND VPWR VPWR _13101_/Y sky130_fd_sc_hd__nand2_1
X_10313_ _10313_/A VGND VGND VPWR VPWR _10313_/Y sky130_fd_sc_hd__inv_2
X_14081_ _14047_/X _14080_/X _14047_/A _14080_/X VGND VGND VPWR VPWR _14082_/B sky130_fd_sc_hd__a2bb2o_1
X_11293_ _11590_/A _11293_/B VGND VGND VPWR VPWR _12362_/A sky130_fd_sc_hd__or2_2
XFILLER_3_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13032_ _14749_/A _13032_/B VGND VGND VPWR VPWR _13032_/X sky130_fd_sc_hd__or2_1
X_10244_ _10244_/A _10244_/B VGND VGND VPWR VPWR _10244_/X sky130_fd_sc_hd__or2_1
XFILLER_105_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10175_ _10175_/A VGND VGND VPWR VPWR _10175_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14983_ _14931_/X _14982_/Y _14964_/Y VGND VGND VPWR VPWR _14983_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13934_ _14644_/A _13838_/B _13838_/Y VGND VGND VPWR VPWR _13934_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13865_ _15113_/A _13865_/B VGND VGND VPWR VPWR _13865_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15604_ _16042_/A VGND VGND VPWR VPWR _15679_/A sky130_fd_sc_hd__inv_2
XFILLER_62_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12816_ _12844_/A _12844_/B VGND VGND VPWR VPWR _12816_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13796_ _13797_/A _13797_/B VGND VGND VPWR VPWR _13798_/A sky130_fd_sc_hd__and2_1
XFILLER_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15535_ _15531_/Y _15616_/A _15534_/Y VGND VGND VPWR VPWR _15540_/B sky130_fd_sc_hd__o21ai_2
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12771_/A _12771_/B VGND VGND VPWR VPWR _12747_/Y sky130_fd_sc_hd__nor2_1
X_15466_ _15399_/X _15465_/X _15399_/X _15465_/X VGND VGND VPWR VPWR _15467_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _11611_/X _12677_/X _11611_/X _12677_/X VGND VGND VPWR VPWR _12679_/B sky130_fd_sc_hd__o2bb2a_1
X_11629_ _11629_/A _11629_/B VGND VGND VPWR VPWR _11629_/Y sky130_fd_sc_hd__nor2_1
X_14417_ _15030_/A _11739_/Y _11777_/Y _14416_/Y VGND VGND VPWR VPWR _14417_/X sky130_fd_sc_hd__o22a_1
X_15397_ _13936_/A _13936_/B _15395_/X _15471_/A VGND VGND VPWR VPWR _15397_/X sky130_fd_sc_hd__a31o_1
X_14348_ _14382_/A _15952_/A VGND VGND VPWR VPWR _15636_/A sky130_fd_sc_hd__and2_1
XFILLER_7_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14279_ _14180_/Y _14277_/Y _14278_/Y VGND VGND VPWR VPWR _14286_/A sky130_fd_sc_hd__o21ai_1
XFILLER_131_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16018_ _15951_/X _16017_/X _15951_/X _16017_/X VGND VGND VPWR VPWR _16034_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08839_/Y _08723_/X _08839_/Y _08723_/X VGND VGND VPWR VPWR _08944_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _09333_/A VGND VGND VPWR VPWR _09486_/A sky130_fd_sc_hd__buf_1
XFILLER_38_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09323_ _09323_/A VGND VGND VPWR VPWR _09328_/A sky130_fd_sc_hd__inv_2
X_09254_ _08916_/A _10102_/B _08935_/X _08935_/A _08935_/B VGND VGND VPWR VPWR _09301_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09185_ _09430_/A _09185_/B VGND VGND VPWR VPWR _09185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08969_ _08965_/Y _11393_/A _08968_/Y VGND VGND VPWR VPWR _08969_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11980_ _11978_/Y _11979_/Y _11936_/Y VGND VGND VPWR VPWR _12069_/A sky130_fd_sc_hd__o21ai_1
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10931_ _09990_/A _09660_/B _09660_/Y VGND VGND VPWR VPWR _10931_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13650_ _13649_/A _13649_/B _13709_/A VGND VGND VPWR VPWR _13650_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10862_ _10438_/A _10861_/A _10438_/Y _10861_/Y _10926_/A VGND VGND VPWR VPWR _12057_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _15512_/A _12322_/B _12322_/X VGND VGND VPWR VPWR _12602_/A sky130_fd_sc_hd__o21ba_1
X_13581_ _12850_/A _13548_/B _13549_/Y _13580_/X VGND VGND VPWR VPWR _13581_/X sky130_fd_sc_hd__o22a_1
X_10793_ _09909_/Y _10791_/X _09911_/A _09910_/Y _10792_/X VGND VGND VPWR VPWR _12938_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ _13440_/A _12309_/B _12309_/Y VGND VGND VPWR VPWR _12533_/B sky130_fd_sc_hd__o21a_1
X_15320_ _15335_/A _15335_/B VGND VGND VPWR VPWR _15384_/A sky130_fd_sc_hd__and2_1
XFILLER_12_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15251_ _15222_/X _15250_/Y _15222_/X _15250_/Y VGND VGND VPWR VPWR _15252_/B sky130_fd_sc_hd__a2bb2o_1
X_12463_ _12459_/X _12462_/X _12459_/X _12462_/X VGND VGND VPWR VPWR _12466_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14202_ _14202_/A _12627_/X VGND VGND VPWR VPWR _14202_/X sky130_fd_sc_hd__or2b_1
X_11414_ _11411_/A _11411_/B _11245_/X _11413_/X VGND VGND VPWR VPWR _13350_/A sky130_fd_sc_hd__o211a_1
XFILLER_125_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12394_ _12393_/A _12458_/B _12393_/Y VGND VGND VPWR VPWR _12394_/X sky130_fd_sc_hd__o21a_1
X_15182_ _15116_/A _15116_/B _15116_/Y VGND VGND VPWR VPWR _15182_/Y sky130_fd_sc_hd__o21ai_1
X_14133_ _14133_/A VGND VGND VPWR VPWR _14133_/Y sky130_fd_sc_hd__inv_2
X_11345_ _13042_/A _11344_/B _11344_/Y VGND VGND VPWR VPWR _11345_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14064_ _14064_/A _14064_/B VGND VGND VPWR VPWR _14064_/X sky130_fd_sc_hd__or2_1
X_11276_ _11276_/A _11276_/B VGND VGND VPWR VPWR _11276_/X sky130_fd_sc_hd__and2_1
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13015_ _13015_/A VGND VGND VPWR VPWR _14493_/A sky130_fd_sc_hd__buf_1
X_10227_ _10309_/B _10226_/X _10309_/B _10226_/X VGND VGND VPWR VPWR _10296_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10158_ _09249_/B _10128_/B _10129_/B VGND VGND VPWR VPWR _10159_/B sky130_fd_sc_hd__a21bo_1
X_14966_ _14931_/X _14965_/Y _14931_/X _14965_/Y VGND VGND VPWR VPWR _14984_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10089_ _09749_/X _10034_/B _10034_/Y _10088_/X VGND VGND VPWR VPWR _10089_/X sky130_fd_sc_hd__a2bb2o_1
X_13917_ _15406_/A _13948_/B VGND VGND VPWR VPWR _13917_/Y sky130_fd_sc_hd__nor2_1
X_14897_ _14817_/X _14896_/X _14817_/X _14896_/X VGND VGND VPWR VPWR _14908_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13848_ _14623_/A _13848_/B VGND VGND VPWR VPWR _13848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13779_ _15116_/A _13779_/B VGND VGND VPWR VPWR _13779_/Y sky130_fd_sc_hd__nor2_1
X_15518_ _15475_/X _15517_/Y _15475_/X _15517_/Y VGND VGND VPWR VPWR _15640_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15449_ _15449_/A _15449_/B VGND VGND VPWR VPWR _15449_/X sky130_fd_sc_hd__and2_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09941_ _09941_/A VGND VGND VPWR VPWR _10792_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09872_ _09448_/Y _09871_/X _09478_/X VGND VGND VPWR VPWR _09873_/A sky130_fd_sc_hd__o21ai_2
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08823_/A VGND VGND VPWR VPWR _08823_/X sky130_fd_sc_hd__buf_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _09331_/A VGND VGND VPWR VPWR _09482_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _09551_/A _08596_/A _08598_/Y _08684_/X VGND VGND VPWR VPWR _08685_/X sky130_fd_sc_hd__o22a_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09306_ _10245_/A _09307_/B VGND VGND VPWR VPWR _09306_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09237_ _08721_/B _09799_/A _09231_/Y _09628_/A VGND VGND VPWR VPWR _09238_/A sky130_fd_sc_hd__o22a_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09168_ _10008_/B _09167_/B _09167_/Y VGND VGND VPWR VPWR _09169_/A sky130_fd_sc_hd__a21oi_2
XFILLER_119_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09099_ _09069_/A _09069_/B _09070_/B VGND VGND VPWR VPWR _09709_/A sky130_fd_sc_hd__o21a_1
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11130_ _12078_/A _11130_/B VGND VGND VPWR VPWR _11130_/X sky130_fd_sc_hd__and2_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11061_ _11061_/A _13754_/B VGND VGND VPWR VPWR _11062_/A sky130_fd_sc_hd__or2_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10012_ _10012_/A _10012_/B VGND VGND VPWR VPWR _10044_/B sky130_fd_sc_hd__nor2_1
X_14820_ _14802_/A _14802_/B _14802_/X _14819_/X VGND VGND VPWR VPWR _14820_/X sky130_fd_sc_hd__o22a_1
XFILLER_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11963_ _13101_/A _11962_/B _11064_/B _11962_/X VGND VGND VPWR VPWR _11963_/X sky130_fd_sc_hd__o22a_1
X_14751_ _14674_/A _14674_/B _14671_/X _14674_/Y VGND VGND VPWR VPWR _14751_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_57_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10914_ _14623_/A _10867_/B _10867_/X _10913_/X VGND VGND VPWR VPWR _10914_/X sky130_fd_sc_hd__o22a_1
XFILLER_72_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14682_ _14682_/A _14681_/X VGND VGND VPWR VPWR _14682_/X sky130_fd_sc_hd__or2b_1
XFILLER_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11894_ _11894_/A VGND VGND VPWR VPWR _11894_/Y sky130_fd_sc_hd__inv_2
X_13702_ _13727_/A _13700_/X _13701_/X VGND VGND VPWR VPWR _13702_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16421_ _16465_/Q VGND VGND VPWR VPWR _16421_/Y sky130_fd_sc_hd__inv_2
X_10845_ _10921_/A _10922_/B VGND VGND VPWR VPWR _11011_/A sky130_fd_sc_hd__and2_1
XFILLER_71_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13633_ _13633_/A VGND VGND VPWR VPWR _15128_/A sky130_fd_sc_hd__buf_1
XFILLER_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16352_ _16333_/X _16351_/Y _16333_/X _16351_/Y VGND VGND VPWR VPWR _16402_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15303_ _14588_/A _15246_/B _15246_/Y VGND VGND VPWR VPWR _15303_/Y sky130_fd_sc_hd__o21ai_1
X_10776_ _13063_/A _10704_/B _10704_/Y _10775_/X VGND VGND VPWR VPWR _10776_/X sky130_fd_sc_hd__a2bb2o_1
X_13564_ _13564_/A _13564_/B VGND VGND VPWR VPWR _13565_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16283_ _16269_/X _16282_/Y _16269_/X _16282_/Y VGND VGND VPWR VPWR _16336_/B sky130_fd_sc_hd__o2bb2a_1
X_12515_ _12514_/A _12514_/B _12514_/Y _11707_/X VGND VGND VPWR VPWR _12635_/A sky130_fd_sc_hd__o211a_1
X_13495_ _13495_/A _13495_/B VGND VGND VPWR VPWR _13495_/X sky130_fd_sc_hd__and2_1
X_15234_ _15234_/A _15234_/B VGND VGND VPWR VPWR _15234_/Y sky130_fd_sc_hd__nand2_1
X_12446_ _12441_/X _12445_/X _12441_/X _12445_/X VGND VGND VPWR VPWR _12447_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15165_ _15100_/X _15105_/A _15104_/X VGND VGND VPWR VPWR _15165_/Y sky130_fd_sc_hd__o21ai_1
X_12377_ _11530_/Y _12376_/X _11530_/Y _12376_/X VGND VGND VPWR VPWR _12379_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14116_ _14079_/Y _14113_/X _14880_/A _14115_/Y VGND VGND VPWR VPWR _14116_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11328_ _09377_/B _10239_/B _10239_/X VGND VGND VPWR VPWR _11329_/B sky130_fd_sc_hd__a21boi_1
XFILLER_99_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15096_ _15063_/A _15063_/B _15063_/Y _15095_/X VGND VGND VPWR VPWR _15096_/X sky130_fd_sc_hd__a2bb2o_1
X_14047_ _14047_/A VGND VGND VPWR VPWR _14047_/X sky130_fd_sc_hd__buf_1
X_11259_ _15449_/A _11197_/B _11197_/Y _11258_/X VGND VGND VPWR VPWR _11259_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15998_ _16053_/A _16053_/B VGND VGND VPWR VPWR _15998_/X sky130_fd_sc_hd__and2_1
XFILLER_67_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14949_ _14949_/A _14948_/X VGND VGND VPWR VPWR _14949_/X sky130_fd_sc_hd__or2b_1
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08470_ input5/X input21/X VGND VGND VPWR VPWR _08470_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09022_ _08795_/X _09011_/Y _08592_/Y _09011_/Y VGND VGND VPWR VPWR _09551_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09924_ _09924_/A VGND VGND VPWR VPWR _09924_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09855_ _09855_/A _09855_/B VGND VGND VPWR VPWR _09855_/X sky130_fd_sc_hd__or2_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08806_ _08806_/A VGND VGND VPWR VPWR _08806_/Y sky130_fd_sc_hd__inv_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09786_ _09995_/B _09784_/Y _09785_/Y VGND VGND VPWR VPWR _09788_/B sky130_fd_sc_hd__o21ai_1
X_08737_ _10011_/A _09529_/A VGND VGND VPWR VPWR _08737_/X sky130_fd_sc_hd__or2_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08668_ _08394_/B _08665_/A _08671_/A _08667_/Y VGND VGND VPWR VPWR _09541_/B sky130_fd_sc_hd__o22a_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10630_ _10612_/Y _10627_/X _10629_/Y VGND VGND VPWR VPWR _10631_/A sky130_fd_sc_hd__o21ai_1
X_08599_ _08599_/A VGND VGND VPWR VPWR _08599_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10561_ _10561_/A VGND VGND VPWR VPWR _10561_/Y sky130_fd_sc_hd__inv_2
X_12300_ _12300_/A _12300_/B VGND VGND VPWR VPWR _12300_/Y sky130_fd_sc_hd__nand2_1
X_13280_ _13260_/Y _13278_/Y _13279_/Y VGND VGND VPWR VPWR _13281_/A sky130_fd_sc_hd__o21ai_2
X_10492_ _10490_/Y _10491_/Y _10491_/A _09846_/X _09941_/A VGND VGND VPWR VPWR _12928_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12231_ _14048_/A VGND VGND VPWR VPWR _13351_/A sky130_fd_sc_hd__inv_2
XFILLER_6_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12162_ _12160_/Y _12161_/Y _12098_/Y VGND VGND VPWR VPWR _12255_/A sky130_fd_sc_hd__o21ai_1
XFILLER_123_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12093_ _09396_/A _12165_/B _09396_/A _12165_/B VGND VGND VPWR VPWR _12093_/X sky130_fd_sc_hd__a2bb2o_1
X_11113_ _11587_/A _11113_/B VGND VGND VPWR VPWR _12252_/A sky130_fd_sc_hd__or2_1
X_15921_ _15964_/A _15964_/B VGND VGND VPWR VPWR _15999_/A sky130_fd_sc_hd__and2_1
XFILLER_110_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11044_ _10883_/A _10883_/B _10883_/A _10883_/B VGND VGND VPWR VPWR _11044_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15852_ _14171_/A _15851_/X _12639_/X VGND VGND VPWR VPWR _15853_/A sky130_fd_sc_hd__o21ai_1
XFILLER_91_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15783_ _16245_/A _16241_/A _15782_/X VGND VGND VPWR VPWR _15788_/B sky130_fd_sc_hd__o21ai_1
X_14803_ _15464_/A VGND VGND VPWR VPWR _14806_/A sky130_fd_sc_hd__buf_1
XFILLER_76_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12995_ _14461_/A _12926_/B _12926_/Y VGND VGND VPWR VPWR _12995_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14734_ _14792_/A _14732_/X _14733_/X VGND VGND VPWR VPWR _14734_/X sky130_fd_sc_hd__o21a_1
X_11946_ _13693_/A _11901_/B _11901_/Y VGND VGND VPWR VPWR _11946_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16404_ _16454_/A _16404_/B VGND VGND VPWR VPWR _16473_/D sky130_fd_sc_hd__or2_1
X_14665_ _14665_/A _14665_/B VGND VGND VPWR VPWR _14665_/Y sky130_fd_sc_hd__nor2_1
X_11877_ _13621_/A _11839_/B _11839_/Y VGND VGND VPWR VPWR _11877_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13616_ _13616_/A VGND VGND VPWR VPWR _13616_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14596_ _12091_/Y _14595_/X _12091_/Y _14595_/X VGND VGND VPWR VPWR _14597_/B sky130_fd_sc_hd__o2bb2a_1
X_10828_ _12080_/A VGND VGND VPWR VPWR _12690_/A sky130_fd_sc_hd__buf_1
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16335_ _16287_/Y _16333_/X _16334_/Y VGND VGND VPWR VPWR _16335_/X sky130_fd_sc_hd__o21a_1
X_10759_ _10764_/A _10758_/X _10764_/A _10758_/X VGND VGND VPWR VPWR _10766_/B sky130_fd_sc_hd__a2bb2o_1
X_13547_ _13537_/X _13546_/Y _13537_/X _13546_/Y VGND VGND VPWR VPWR _13548_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16266_ _16266_/A _16266_/B VGND VGND VPWR VPWR _16266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13478_ _14309_/A _13478_/B VGND VGND VPWR VPWR _15982_/A sky130_fd_sc_hd__or2_1
X_15217_ _15212_/X _15268_/A _15216_/X VGND VGND VPWR VPWR _15217_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16197_ _16197_/A VGND VGND VPWR VPWR _16197_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12429_ _12429_/A VGND VGND VPWR VPWR _12429_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15148_ _15143_/A _15143_/B _15143_/Y _15147_/X VGND VGND VPWR VPWR _15148_/X sky130_fd_sc_hd__a2bb2o_1
X_15079_ _15079_/A _15030_/X VGND VGND VPWR VPWR _15079_/X sky130_fd_sc_hd__or2b_1
XFILLER_68_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09640_ _09958_/A _09640_/B VGND VGND VPWR VPWR _09640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09571_ _09516_/X _09570_/X _09516_/X _09570_/X VGND VGND VPWR VPWR _09997_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_82_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08522_ _09862_/A VGND VGND VPWR VPWR _09348_/B sky130_fd_sc_hd__inv_2
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08453_ _08453_/A VGND VGND VPWR VPWR _08453_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08384_ _08384_/A VGND VGND VPWR VPWR _08384_/Y sky130_fd_sc_hd__inv_2
X_09005_ _08935_/A _09232_/B _08664_/X VGND VGND VPWR VPWR _09005_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09907_ _10654_/B _09906_/X VGND VGND VPWR VPWR _09908_/B sky130_fd_sc_hd__or2b_1
XFILLER_76_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _09838_/A _09838_/B VGND VGND VPWR VPWR _09839_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09769_ _09769_/A VGND VGND VPWR VPWR _09773_/A sky130_fd_sc_hd__inv_2
X_11800_ _11798_/A _11798_/B _11798_/X _11799_/Y VGND VGND VPWR VPWR _11847_/B sky130_fd_sc_hd__a22o_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12735_/Y _12778_/X _12779_/Y VGND VGND VPWR VPWR _12780_/X sky130_fd_sc_hd__o21a_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11731_ _11731_/A _11731_/B VGND VGND VPWR VPWR _11731_/Y sky130_fd_sc_hd__nor2_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14433_/X _14449_/X _14433_/X _14449_/X VGND VGND VPWR VPWR _14463_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11662_ _09196_/Y _09193_/A _09198_/X _09193_/Y VGND VGND VPWR VPWR _11663_/A sky130_fd_sc_hd__o22a_1
X_14381_ _15644_/A _14379_/X _14380_/X VGND VGND VPWR VPWR _14381_/X sky130_fd_sc_hd__o21a_1
X_13401_ _14091_/A VGND VGND VPWR VPWR _14908_/A sky130_fd_sc_hd__buf_1
X_11593_ _12444_/A VGND VGND VPWR VPWR _12863_/A sky130_fd_sc_hd__inv_2
X_10613_ _08928_/A _10277_/Y _08929_/B _10277_/A VGND VGND VPWR VPWR _10756_/B sky130_fd_sc_hd__o22a_1
X_16120_ _16116_/Y _16147_/A _16119_/Y VGND VGND VPWR VPWR _16140_/A sky130_fd_sc_hd__o21ai_2
X_13332_ _14731_/A _13285_/B _13285_/Y VGND VGND VPWR VPWR _13332_/Y sky130_fd_sc_hd__o21ai_1
X_10544_ _11801_/A _10544_/B VGND VGND VPWR VPWR _10544_/X sky130_fd_sc_hd__and2_1
XFILLER_22_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16051_ _16051_/A _16051_/B VGND VGND VPWR VPWR _16051_/Y sky130_fd_sc_hd__nand2_1
X_13263_ _13185_/X _13262_/Y _13185_/X _13262_/Y VGND VGND VPWR VPWR _13276_/B sky130_fd_sc_hd__a2bb2o_1
X_10475_ _10552_/A _11852_/A VGND VGND VPWR VPWR _10475_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12214_ _12146_/X _12213_/X _12146_/X _12213_/X VGND VGND VPWR VPWR _12215_/B sky130_fd_sc_hd__a2bb2o_1
X_13194_ _13194_/A _13194_/B VGND VGND VPWR VPWR _13194_/Y sky130_fd_sc_hd__nand2_1
X_15002_ _11811_/A _15001_/X _11810_/X VGND VGND VPWR VPWR _15002_/X sky130_fd_sc_hd__o21a_1
X_12145_ _13914_/A _12145_/B VGND VGND VPWR VPWR _12145_/X sky130_fd_sc_hd__or2_1
XFILLER_1_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12076_ _12076_/A VGND VGND VPWR VPWR _12076_/Y sky130_fd_sc_hd__inv_2
X_15904_ _15906_/A _15906_/B VGND VGND VPWR VPWR _15904_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11027_ _13910_/A _11087_/B VGND VGND VPWR VPWR _11210_/A sky130_fd_sc_hd__and2_1
XFILLER_77_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15835_ _15822_/X _15834_/X _15822_/X _15834_/X VGND VGND VPWR VPWR _15836_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15766_ _14906_/A _14906_/B _14906_/Y VGND VGND VPWR VPWR _15766_/X sky130_fd_sc_hd__o21a_1
X_12978_ _13697_/A VGND VGND VPWR VPWR _14481_/A sky130_fd_sc_hd__inv_2
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15697_ _15578_/Y _15695_/X _15696_/Y VGND VGND VPWR VPWR _15697_/X sky130_fd_sc_hd__o21a_1
X_14717_ _14645_/Y _14716_/X _14645_/Y _14716_/X VGND VGND VPWR VPWR _14718_/B sky130_fd_sc_hd__a2bb2o_1
X_11929_ _12775_/A _11986_/A _11928_/Y VGND VGND VPWR VPWR _11929_/Y sky130_fd_sc_hd__a21oi_1
X_14648_ _15333_/A _14648_/B VGND VGND VPWR VPWR _14648_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16318_ _16318_/A _16318_/B VGND VGND VPWR VPWR _16318_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14579_ _14559_/Y _14577_/X _14578_/Y VGND VGND VPWR VPWR _14579_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16249_ _16249_/A _16249_/B VGND VGND VPWR VPWR _16249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09623_ _09506_/X _09622_/X _09506_/X _09622_/X VGND VGND VPWR VPWR _09957_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09554_ _09601_/A _09552_/X _09601_/B VGND VGND VPWR VPWR _09554_/X sky130_fd_sc_hd__o21ba_1
XFILLER_24_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09485_ _08773_/A _09473_/X _08773_/A _09473_/X VGND VGND VPWR VPWR _09486_/B sky130_fd_sc_hd__o2bb2a_1
X_08505_ _09146_/A _08505_/B VGND VGND VPWR VPWR _08508_/A sky130_fd_sc_hd__or2_1
XFILLER_24_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08436_ _10012_/A VGND VGND VPWR VPWR _08712_/A sky130_fd_sc_hd__inv_2
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08367_ _08272_/A input11/X _08364_/B _08366_/A VGND VGND VPWR VPWR _08409_/A sky130_fd_sc_hd__o22a_1
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08298_ _08298_/A VGND VGND VPWR VPWR _08298_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10260_ _09328_/B _10241_/B _10241_/X _10981_/A VGND VGND VPWR VPWR _11155_/A sky130_fd_sc_hd__a22o_1
XFILLER_117_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10191_ _10239_/B _10143_/B _10143_/Y _11322_/A VGND VGND VPWR VPWR _10191_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_120_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13950_ _15408_/A _13950_/B VGND VGND VPWR VPWR _13950_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12901_ _12842_/A _12842_/B _12842_/Y VGND VGND VPWR VPWR _12901_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _15620_/A _14386_/X VGND VGND VPWR VPWR _15620_/X sky130_fd_sc_hd__or2b_1
X_13881_ _13863_/X _13880_/Y _13863_/X _13880_/Y VGND VGND VPWR VPWR _13883_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12832_ _12832_/A _12832_/B VGND VGND VPWR VPWR _12832_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15494_/X _15549_/X _15690_/B VGND VGND VPWR VPWR _15551_/X sky130_fd_sc_hd__o21a_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12763_/A _12763_/B VGND VGND VPWR VPWR _12763_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15482_ _14786_/A _15449_/B _15449_/X _15481_/X VGND VGND VPWR VPWR _15482_/X sky130_fd_sc_hd__o22a_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14459_/A _14459_/B _14459_/Y VGND VGND VPWR VPWR _14502_/X sky130_fd_sc_hd__o21a_1
X_11714_ _11713_/A _11720_/B _11713_/Y VGND VGND VPWR VPWR _11716_/A sky130_fd_sc_hd__a21oi_2
XFILLER_30_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14427_/A _14427_/B _14427_/X _14432_/X VGND VGND VPWR VPWR _14433_/X sky130_fd_sc_hd__o22a_1
XFILLER_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12694_ _12694_/A _12694_/B VGND VGND VPWR VPWR _12694_/Y sky130_fd_sc_hd__nor2_1
X_11645_ _11642_/X _11644_/Y _11642_/X _11644_/Y VGND VGND VPWR VPWR _11647_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 wbs_adr_i[7] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_4
XFILLER_128_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14364_ _14364_/A _15774_/A VGND VGND VPWR VPWR _14376_/A sky130_fd_sc_hd__or2_1
X_11576_ _11576_/A _11576_/B VGND VGND VPWR VPWR _11576_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput26 wbs_dat_i[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_4
X_16103_ _16035_/X _16102_/Y _16035_/X _16102_/Y VGND VGND VPWR VPWR _16103_/X sky130_fd_sc_hd__a2bb2o_1
X_14295_ _14295_/A _14288_/X VGND VGND VPWR VPWR _14295_/X sky130_fd_sc_hd__or2b_1
X_13315_ _13302_/A _13314_/Y _13302_/A _13314_/Y VGND VGND VPWR VPWR _13371_/B sky130_fd_sc_hd__a2bb2o_1
X_10527_ _11837_/A _10527_/B VGND VGND VPWR VPWR _10527_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16034_ _16034_/A _16034_/B VGND VGND VPWR VPWR _16034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13246_ _15072_/A VGND VGND VPWR VPWR _14421_/A sky130_fd_sc_hd__inv_2
X_10458_ _10966_/A _11213_/A VGND VGND VPWR VPWR _10459_/A sky130_fd_sc_hd__or2_1
XFILLER_111_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13177_ _13102_/X _13176_/Y _13102_/X _13176_/Y VGND VGND VPWR VPWR _13184_/B sky130_fd_sc_hd__a2bb2o_1
X_10389_ _10368_/X _10388_/X _10368_/X _10388_/X VGND VGND VPWR VPWR _10442_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12128_ _15081_/A _12139_/B VGND VGND VPWR VPWR _12225_/A sky130_fd_sc_hd__and2_1
XFILLER_111_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12059_ _12059_/A _12059_/B VGND VGND VPWR VPWR _12059_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15818_ _15725_/Y _15816_/X _15817_/Y VGND VGND VPWR VPWR _15818_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15749_ _16108_/A _15809_/B VGND VGND VPWR VPWR _15749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09270_ _08597_/A _09856_/A _09216_/A VGND VGND VPWR VPWR _09270_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ _08875_/X _08983_/X _11460_/B VGND VGND VPWR VPWR _08985_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09606_ _09980_/A VGND VGND VPWR VPWR _09981_/A sky130_fd_sc_hd__buf_1
XFILLER_71_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09537_ _09547_/A _09547_/B VGND VGND VPWR VPWR _09648_/A sky130_fd_sc_hd__nor2_1
XFILLER_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09468_ _09454_/Y _09466_/X _09467_/X VGND VGND VPWR VPWR _09468_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09399_ _15060_/A VGND VGND VPWR VPWR _13898_/A sky130_fd_sc_hd__buf_1
XFILLER_8_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08419_ _08419_/A VGND VGND VPWR VPWR _08441_/A sky130_fd_sc_hd__clkbuf_2
X_11430_ _12586_/A _12585_/A _11429_/X VGND VGND VPWR VPWR _11434_/B sky130_fd_sc_hd__o21ai_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11361_ _14062_/A _11179_/B _11179_/Y VGND VGND VPWR VPWR _11361_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13100_ _14568_/A _13101_/B VGND VGND VPWR VPWR _13100_/Y sky130_fd_sc_hd__nor2_1
X_10312_ _10247_/A _10247_/B _10247_/X VGND VGND VPWR VPWR _10313_/A sky130_fd_sc_hd__o21ba_1
XFILLER_106_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14080_ _14815_/A _14048_/B _14048_/Y VGND VGND VPWR VPWR _14080_/X sky130_fd_sc_hd__a21o_1
X_11292_ _09995_/B _11291_/X _09995_/B _11291_/X VGND VGND VPWR VPWR _11293_/B sky130_fd_sc_hd__a2bb2o_1
X_13031_ _13050_/A _13029_/X _13030_/X VGND VGND VPWR VPWR _13031_/X sky130_fd_sc_hd__o21a_1
X_10243_ _10243_/A _10243_/B VGND VGND VPWR VPWR _10243_/X sky130_fd_sc_hd__or2_1
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10174_ _10100_/Y _08647_/A _10111_/A VGND VGND VPWR VPWR _10175_/A sky130_fd_sc_hd__o21ai_2
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14982_ _15563_/A _14982_/B VGND VGND VPWR VPWR _14982_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13933_ _14430_/A VGND VGND VPWR VPWR _15396_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13864_ _13864_/A VGND VGND VPWR VPWR _13864_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15603_ _15602_/A _15601_/Y _15602_/Y _15601_/A _15595_/A VGND VGND VPWR VPWR _16042_/A
+ sky130_fd_sc_hd__a221o_1
X_12815_ _12768_/X _12814_/Y _12768_/X _12814_/Y VGND VGND VPWR VPWR _12844_/B sky130_fd_sc_hd__a2bb2o_1
X_15534_ _15534_/A _15534_/B VGND VGND VPWR VPWR _15534_/Y sky130_fd_sc_hd__nand2_1
X_13795_ _13777_/X _13794_/X _13777_/X _13794_/X VGND VGND VPWR VPWR _13797_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12712_/X _12745_/X _12712_/X _12745_/X VGND VGND VPWR VPWR _12771_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15465_ _15465_/A _15400_/X VGND VGND VPWR VPWR _15465_/X sky130_fd_sc_hd__or2b_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _11612_/Y _12676_/Y _11528_/X VGND VGND VPWR VPWR _12677_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15396_ _15396_/A _15396_/B VGND VGND VPWR VPWR _15471_/A sky130_fd_sc_hd__and2_1
X_14416_ _14416_/A VGND VGND VPWR VPWR _14416_/Y sky130_fd_sc_hd__inv_2
X_11628_ _11625_/Y _11627_/X _11625_/Y _11627_/X VGND VGND VPWR VPWR _11629_/B sky130_fd_sc_hd__o2bb2a_1
X_14347_ _14353_/A _14347_/B VGND VGND VPWR VPWR _15952_/A sky130_fd_sc_hd__or2_1
XFILLER_7_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11559_ _11559_/A _11558_/X VGND VGND VPWR VPWR _11559_/X sky130_fd_sc_hd__or2b_1
XFILLER_116_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14278_ _14278_/A _14278_/B VGND VGND VPWR VPWR _14278_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16017_ _16017_/A _15952_/X VGND VGND VPWR VPWR _16017_/X sky130_fd_sc_hd__or2b_1
X_13229_ _13199_/X _13228_/Y _13199_/X _13228_/Y VGND VGND VPWR VPWR _13297_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _08770_/A _08770_/B VGND VGND VPWR VPWR _08770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09322_ _09319_/X _09321_/X _09319_/X _09321_/X VGND VGND VPWR VPWR _09323_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09253_ _09458_/A _09253_/B VGND VGND VPWR VPWR _10061_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09184_ _09184_/A VGND VGND VPWR VPWR _09184_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08968_ _08968_/A _08968_/B VGND VGND VPWR VPWR _08968_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08899_ _10014_/A _09249_/B _08803_/Y VGND VGND VPWR VPWR _08899_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10930_ _10930_/A VGND VGND VPWR VPWR _11587_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12600_ _12600_/A VGND VGND VPWR VPWR _12600_/Y sky130_fd_sc_hd__inv_2
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10861_ _10861_/A VGND VGND VPWR VPWR _10861_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13580_ _12848_/A _13552_/B _13553_/Y _13579_/X VGND VGND VPWR VPWR _13580_/X sky130_fd_sc_hd__o22a_1
X_10792_ _10792_/A VGND VGND VPWR VPWR _10792_/X sky130_fd_sc_hd__clkbuf_2
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ _12530_/A _12530_/B _12530_/Y _11707_/A VGND VGND VPWR VPWR _12631_/A sky130_fd_sc_hd__o211a_1
XFILLER_12_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15250_ _15196_/A _15196_/B _15196_/Y VGND VGND VPWR VPWR _15250_/Y sky130_fd_sc_hd__o21ai_1
X_12462_ _12462_/A _12460_/X VGND VGND VPWR VPWR _12462_/X sky130_fd_sc_hd__or2b_1
X_14201_ _14207_/A _14201_/B VGND VGND VPWR VPWR _15866_/A sky130_fd_sc_hd__or2_1
X_11413_ _13936_/A _12232_/B VGND VGND VPWR VPWR _11413_/X sky130_fd_sc_hd__or2_1
X_15181_ _15181_/A _15181_/B VGND VGND VPWR VPWR _15181_/Y sky130_fd_sc_hd__nand2_1
X_12393_ _12393_/A _12458_/B VGND VGND VPWR VPWR _12393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14132_ _14132_/A VGND VGND VPWR VPWR _14868_/A sky130_fd_sc_hd__inv_2
X_11344_ _13042_/A _11344_/B VGND VGND VPWR VPWR _11344_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14063_ _14129_/A _14061_/X _14062_/X VGND VGND VPWR VPWR _14063_/X sky130_fd_sc_hd__o21a_1
X_11275_ _15054_/A VGND VGND VPWR VPWR _13890_/A sky130_fd_sc_hd__buf_1
XFILLER_79_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13014_ _13090_/A _13011_/X _13013_/X VGND VGND VPWR VPWR _13014_/X sky130_fd_sc_hd__o21a_1
X_10226_ _10226_/A VGND VGND VPWR VPWR _10226_/X sky130_fd_sc_hd__buf_1
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10157_ _10159_/A VGND VGND VPWR VPWR _10243_/B sky130_fd_sc_hd__buf_1
X_14965_ _15563_/A _14982_/B _14964_/Y VGND VGND VPWR VPWR _14965_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_82_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10088_ _10037_/X _10086_/X _11520_/B VGND VGND VPWR VPWR _10088_/X sky130_fd_sc_hd__o21a_1
X_13916_ _13847_/X _13915_/Y _13847_/X _13915_/Y VGND VGND VPWR VPWR _13948_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14896_ _14809_/A _14809_/B _14809_/Y VGND VGND VPWR VPWR _14896_/X sky130_fd_sc_hd__a21o_1
XFILLER_75_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13847_ _13821_/Y _13845_/X _13846_/Y VGND VGND VPWR VPWR _13847_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13778_ _13778_/A VGND VGND VPWR VPWR _13778_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15517_ _15467_/A _15467_/B _15467_/Y VGND VGND VPWR VPWR _15517_/Y sky130_fd_sc_hd__o21ai_1
X_12729_ _12783_/A _12783_/B VGND VGND VPWR VPWR _12729_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15448_ _15411_/X _15447_/X _15411_/X _15447_/X VGND VGND VPWR VPWR _15449_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15379_ _15338_/X _15378_/X _15338_/X _15378_/X VGND VGND VPWR VPWR _15406_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09940_ _11592_/A VGND VGND VPWR VPWR _09941_/A sky130_fd_sc_hd__inv_2
XFILLER_97_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09871_ _09449_/Y _09870_/X _09476_/X VGND VGND VPWR VPWR _09871_/X sky130_fd_sc_hd__o21a_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _08822_/A VGND VGND VPWR VPWR _08823_/A sky130_fd_sc_hd__inv_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _09478_/A _10134_/A _08752_/X VGND VGND VPWR VPWR _08753_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08684_ _09549_/A _08609_/A _08611_/Y _08683_/X VGND VGND VPWR VPWR _08684_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09305_ _10402_/A _09303_/Y _09304_/Y VGND VGND VPWR VPWR _09307_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09236_ _09629_/A VGND VGND VPWR VPWR _09628_/A sky130_fd_sc_hd__inv_2
XFILLER_119_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09167_ _10008_/B _09167_/B VGND VGND VPWR VPWR _09167_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09098_ _09409_/A VGND VGND VPWR VPWR _09714_/A sky130_fd_sc_hd__inv_2
XFILLER_122_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11060_ _11063_/B VGND VGND VPWR VPWR _13754_/B sky130_fd_sc_hd__inv_2
XFILLER_1_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10011_ _10011_/A _10011_/B VGND VGND VPWR VPWR _10041_/B sky130_fd_sc_hd__nor2_1
XFILLER_130_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14750_ _14677_/A _14677_/B _14670_/X _14677_/Y VGND VGND VPWR VPWR _14750_/X sky130_fd_sc_hd__o2bb2a_1
X_11962_ _13101_/A _11962_/B VGND VGND VPWR VPWR _11962_/X sky130_fd_sc_hd__and2_1
X_13701_ _13701_/A _13701_/B VGND VGND VPWR VPWR _13701_/X sky130_fd_sc_hd__or2_1
XFILLER_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10913_ _14627_/A _10875_/B _10875_/X _10912_/X VGND VGND VPWR VPWR _10913_/X sky130_fd_sc_hd__o22a_1
X_14681_ _15184_/A _14681_/B VGND VGND VPWR VPWR _14681_/X sky130_fd_sc_hd__or2_1
X_11893_ _11885_/Y _11891_/X _11892_/Y VGND VGND VPWR VPWR _11894_/A sky130_fd_sc_hd__o21ai_1
XFILLER_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16420_ _16437_/B _16429_/B VGND VGND VPWR VPWR _16420_/X sky130_fd_sc_hd__or2_1
XFILLER_72_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10844_ _10776_/X _10843_/Y _10776_/X _10843_/Y VGND VGND VPWR VPWR _10922_/B sky130_fd_sc_hd__o2bb2a_1
X_13632_ _13632_/A VGND VGND VPWR VPWR _13632_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16351_ _16334_/A _16334_/B _16334_/Y VGND VGND VPWR VPWR _16351_/Y sky130_fd_sc_hd__o21ai_1
X_13563_ _13533_/X _13562_/Y _13533_/X _13562_/Y VGND VGND VPWR VPWR _13564_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12514_ _12514_/A _12514_/B VGND VGND VPWR VPWR _12514_/Y sky130_fd_sc_hd__nand2_1
X_15302_ _15347_/A _15347_/B VGND VGND VPWR VPWR _15366_/A sky130_fd_sc_hd__and2_1
X_10775_ _13068_/A _10712_/B _10712_/Y _10774_/X VGND VGND VPWR VPWR _10775_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16282_ _16270_/A _16336_/A _16270_/Y VGND VGND VPWR VPWR _16282_/Y sky130_fd_sc_hd__o21ai_1
X_13494_ _11617_/Y _13493_/X _11617_/Y _13493_/X VGND VGND VPWR VPWR _13495_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15233_ _15228_/X _15232_/Y _15228_/X _15232_/Y VGND VGND VPWR VPWR _15234_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12445_ _13133_/A _12439_/B _13133_/A _12439_/B VGND VGND VPWR VPWR _12445_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15164_ _12428_/A _15163_/B _15163_/Y VGND VGND VPWR VPWR _15164_/X sky130_fd_sc_hd__a21o_1
X_12376_ _11518_/A _12270_/Y _12375_/Y VGND VGND VPWR VPWR _12376_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14115_ _14115_/A VGND VGND VPWR VPWR _14115_/Y sky130_fd_sc_hd__inv_2
X_11327_ _11315_/X _11326_/Y _11315_/X _11326_/Y VGND VGND VPWR VPWR _11516_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_125_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15095_ _15066_/A _15066_/B _15066_/Y _15094_/X VGND VGND VPWR VPWR _15095_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11258_ _15452_/A _11206_/B _11206_/Y _11257_/X VGND VGND VPWR VPWR _11258_/X sky130_fd_sc_hd__a2bb2o_1
X_14046_ _13937_/X _14045_/X _13937_/A _14045_/X VGND VGND VPWR VPWR _14048_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10209_ _10903_/A _10215_/A VGND VGND VPWR VPWR _10210_/A sky130_fd_sc_hd__or2_1
X_11189_ _09426_/A _09136_/B _09136_/Y VGND VGND VPWR VPWR _11190_/A sky130_fd_sc_hd__o21ai_1
XFILLER_95_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15997_ _15969_/Y _15996_/X _15969_/Y _15996_/X VGND VGND VPWR VPWR _16053_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_82_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14948_ _14948_/A _14948_/B VGND VGND VPWR VPWR _14948_/X sky130_fd_sc_hd__or2_1
X_14879_ _15544_/A _14920_/B VGND VGND VPWR VPWR _14879_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09021_ _08580_/X _08893_/X _09021_/S VGND VGND VPWR VPWR _09553_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09923_ _09923_/A _09923_/B VGND VGND VPWR VPWR _11298_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09854_ _09855_/A _09897_/A VGND VGND VPWR VPWR _09854_/Y sky130_fd_sc_hd__nor2_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08805_ _08794_/A _09467_/B _08714_/Y VGND VGND VPWR VPWR _08806_/A sky130_fd_sc_hd__a21oi_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09785_ _09785_/A _09785_/B VGND VGND VPWR VPWR _09785_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08736_ _08736_/A VGND VGND VPWR VPWR _08736_/Y sky130_fd_sc_hd__inv_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08667_ _08667_/A VGND VGND VPWR VPWR _08667_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08598_ _08598_/A VGND VGND VPWR VPWR _08598_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10560_ _10244_/B _10163_/B _10163_/Y VGND VGND VPWR VPWR _10561_/A sky130_fd_sc_hd__a21oi_1
XFILLER_127_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10491_ _10491_/A _10491_/B VGND VGND VPWR VPWR _10491_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09219_ _09549_/A _09696_/A VGND VGND VPWR VPWR _09220_/A sky130_fd_sc_hd__or2_1
XFILLER_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12230_ _12230_/A _12230_/B VGND VGND VPWR VPWR _12230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12161_ _12161_/A VGND VGND VPWR VPWR _12161_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12092_ _12167_/B _12091_/Y _12167_/B _12091_/Y VGND VGND VPWR VPWR _12165_/B sky130_fd_sc_hd__o2bb2a_1
X_11112_ _09661_/X _11111_/X _09661_/X _11111_/X VGND VGND VPWR VPWR _11113_/B sky130_fd_sc_hd__a2bb2oi_1
X_15920_ _15901_/X _15919_/Y _15901_/X _15919_/Y VGND VGND VPWR VPWR _15964_/B sky130_fd_sc_hd__a2bb2o_1
X_11043_ _15078_/A VGND VGND VPWR VPWR _13922_/A sky130_fd_sc_hd__buf_1
XFILLER_77_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15851_ _14284_/A _15850_/X _12637_/X VGND VGND VPWR VPWR _15851_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14802_ _14802_/A _14802_/B VGND VGND VPWR VPWR _14802_/X sky130_fd_sc_hd__and2_1
XFILLER_77_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15782_ _15782_/A _15782_/B VGND VGND VPWR VPWR _15782_/X sky130_fd_sc_hd__or2_1
XFILLER_92_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12994_ _12994_/A VGND VGND VPWR VPWR _13012_/A sky130_fd_sc_hd__inv_2
XFILLER_57_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14733_ _14733_/A _14733_/B VGND VGND VPWR VPWR _14733_/X sky130_fd_sc_hd__or2_1
X_11945_ _11945_/A _11972_/B VGND VGND VPWR VPWR _11945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14664_ _14664_/A VGND VGND VPWR VPWR _15349_/A sky130_fd_sc_hd__buf_1
XFILLER_45_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16403_ _16393_/Y _16401_/X _16349_/X _16402_/X VGND VGND VPWR VPWR _16404_/B sky130_fd_sc_hd__o31a_1
X_13615_ _10428_/X _13614_/X _10428_/X _13614_/X VGND VGND VPWR VPWR _13616_/A sky130_fd_sc_hd__a2bb2o_1
X_11876_ _11901_/A _11901_/B VGND VGND VPWR VPWR _11876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14595_ _15042_/A _12076_/Y _12000_/Y _14527_/X VGND VGND VPWR VPWR _14595_/X sky130_fd_sc_hd__o22a_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10827_ _10826_/A _10826_/B _10826_/Y _10982_/A VGND VGND VPWR VPWR _12080_/A sky130_fd_sc_hd__o211a_1
X_16334_ _16334_/A _16334_/B VGND VGND VPWR VPWR _16334_/Y sky130_fd_sc_hd__nand2_1
X_10758_ _13001_/A _10626_/B _10626_/Y VGND VGND VPWR VPWR _10758_/X sky130_fd_sc_hd__a21o_1
X_13546_ _15040_/A _13513_/B _13513_/Y VGND VGND VPWR VPWR _13546_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16265_ _16178_/Y _16263_/X _16264_/Y VGND VGND VPWR VPWR _16265_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13477_ _13449_/X _13476_/X _13449_/X _13476_/X VGND VGND VPWR VPWR _13478_/B sky130_fd_sc_hd__a2bb2oi_1
X_15216_ _15216_/A _15216_/B VGND VGND VPWR VPWR _15216_/X sky130_fd_sc_hd__or2_1
X_12428_ _12428_/A _12432_/B VGND VGND VPWR VPWR _12428_/X sky130_fd_sc_hd__or2_1
X_10689_ _10688_/A _10688_/B _10688_/Y _10982_/A VGND VGND VPWR VPWR _11990_/A sky130_fd_sc_hd__o211a_1
X_16196_ _16196_/A VGND VGND VPWR VPWR _16196_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12359_ _12358_/Y _12250_/X _12290_/Y VGND VGND VPWR VPWR _12359_/X sky130_fd_sc_hd__o21a_1
X_15147_ _15146_/A _15146_/B _10522_/Y _15146_/Y VGND VGND VPWR VPWR _15147_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15078_ _15078_/A _15078_/B VGND VGND VPWR VPWR _15078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14029_ _14032_/A VGND VGND VPWR VPWR _15461_/A sky130_fd_sc_hd__buf_1
XFILLER_101_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09570_ _09482_/A _09482_/B _09482_/Y VGND VGND VPWR VPWR _09570_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08521_ _08697_/A _08521_/B VGND VGND VPWR VPWR _09862_/A sky130_fd_sc_hd__or2_2
XFILLER_51_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08452_ _08543_/B _08446_/Y _09332_/A VGND VGND VPWR VPWR _08453_/A sky130_fd_sc_hd__o21ai_1
XFILLER_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08383_ _08642_/A VGND VGND VPWR VPWR _09228_/A sky130_fd_sc_hd__buf_1
X_09004_ _12300_/A VGND VGND VPWR VPWR _14138_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09906_ _10654_/A _10653_/A VGND VGND VPWR VPWR _09906_/X sky130_fd_sc_hd__or2_1
XFILLER_116_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _09832_/A _09832_/B _09833_/Y _09836_/Y VGND VGND VPWR VPWR _09838_/B sky130_fd_sc_hd__o22a_1
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09768_ _10052_/A VGND VGND VPWR VPWR _10077_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08719_ _08944_/A _08719_/B VGND VGND VPWR VPWR _08719_/Y sky130_fd_sc_hd__nor2_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11730_ _11730_/A VGND VGND VPWR VPWR _11730_/Y sky130_fd_sc_hd__inv_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09699_ _09698_/A _09698_/B _09730_/A VGND VGND VPWR VPWR _09700_/A sky130_fd_sc_hd__a21bo_2
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11659_/X _11685_/A _11659_/X _11685_/A VGND VGND VPWR VPWR _11668_/A sky130_fd_sc_hd__o2bb2a_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14380_ _14380_/A _15950_/A VGND VGND VPWR VPWR _14380_/X sky130_fd_sc_hd__or2_1
X_13400_ _15519_/A VGND VGND VPWR VPWR _14091_/A sky130_fd_sc_hd__inv_2
X_10612_ _10628_/A _10629_/B VGND VGND VPWR VPWR _10612_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11592_ _11592_/A _11592_/B VGND VGND VPWR VPWR _12444_/A sky130_fd_sc_hd__or2_2
XFILLER_22_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13331_ _13331_/A _13331_/B VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__and2_1
X_10543_ _11021_/A VGND VGND VPWR VPWR _10543_/X sky130_fd_sc_hd__buf_1
XFILLER_6_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16050_ _15968_/X _16049_/Y _15968_/X _16049_/Y VGND VGND VPWR VPWR _16050_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13262_ _13825_/A _13186_/B _13186_/Y VGND VGND VPWR VPWR _13262_/Y sky130_fd_sc_hd__o21ai_1
X_15001_ _11765_/A _15000_/X _11764_/X VGND VGND VPWR VPWR _15001_/X sky130_fd_sc_hd__o21a_1
X_10474_ _11852_/A VGND VGND VPWR VPWR _12696_/A sky130_fd_sc_hd__buf_1
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12213_ _12213_/A _12147_/X VGND VGND VPWR VPWR _12213_/X sky130_fd_sc_hd__or2b_1
X_13193_ _13165_/Y _13191_/X _13192_/Y VGND VGND VPWR VPWR _13193_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12144_ _12219_/A _12142_/X _12143_/X VGND VGND VPWR VPWR _12144_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12075_ _12075_/A _12075_/B VGND VGND VPWR VPWR _12075_/X sky130_fd_sc_hd__or2_1
X_15903_ _15859_/Y _15901_/X _15902_/Y VGND VGND VPWR VPWR _15906_/B sky130_fd_sc_hd__o21a_1
X_11026_ _10914_/X _11025_/X _10914_/X _11025_/X VGND VGND VPWR VPWR _11087_/B sky130_fd_sc_hd__a2bb2o_1
X_15834_ _15706_/X _15834_/B VGND VGND VPWR VPWR _15834_/X sky130_fd_sc_hd__and2b_1
XFILLER_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15765_ _15765_/A _15765_/B VGND VGND VPWR VPWR _15793_/A sky130_fd_sc_hd__or2_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12977_ _14412_/A _13024_/B VGND VGND VPWR VPWR _13065_/A sky130_fd_sc_hd__and2_1
XFILLER_18_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15696_ _16055_/A _15696_/B VGND VGND VPWR VPWR _15696_/Y sky130_fd_sc_hd__nand2_1
X_14716_ _14716_/A _14646_/X VGND VGND VPWR VPWR _14716_/X sky130_fd_sc_hd__or2b_1
XFILLER_72_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11928_ _12775_/A _11986_/A VGND VGND VPWR VPWR _11928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14647_ _14716_/A _14645_/Y _14646_/X VGND VGND VPWR VPWR _14647_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11859_ _11859_/A _11859_/B VGND VGND VPWR VPWR _11859_/X sky130_fd_sc_hd__or2_1
X_14578_ _14578_/A _14578_/B VGND VGND VPWR VPWR _14578_/Y sky130_fd_sc_hd__nand2_1
X_16317_ _16312_/Y _16315_/Y _16316_/Y VGND VGND VPWR VPWR _16317_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13529_ _10336_/Y _13481_/A _10336_/Y _13481_/A VGND VGND VPWR VPWR _13530_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16248_ _16457_/S _16248_/B VGND VGND VPWR VPWR _16248_/Y sky130_fd_sc_hd__nor2_1
X_16179_ _16076_/X _16179_/B VGND VGND VPWR VPWR _16179_/X sky130_fd_sc_hd__and2b_1
XFILLER_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09622_ _09502_/A _09502_/B _09502_/Y VGND VGND VPWR VPWR _09622_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09553_ _09553_/A _09553_/B VGND VGND VPWR VPWR _09601_/B sky130_fd_sc_hd__and2_1
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08504_ _09448_/B VGND VGND VPWR VPWR _09561_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09484_ _09484_/A _09484_/B VGND VGND VPWR VPWR _09484_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08435_ _08434_/A _08328_/Y _08434_/Y _08328_/A _08441_/A VGND VGND VPWR VPWR _10012_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_24_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08366_ _08366_/A VGND VGND VPWR VPWR _08366_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08297_ input24/X input8/X input24/X input8/X VGND VGND VPWR VPWR _08298_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10190_ _10240_/B _10147_/B _10147_/Y _11148_/A VGND VGND VPWR VPWR _11322_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_127_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13880_ _14836_/A _13981_/B _13879_/Y VGND VGND VPWR VPWR _13880_/Y sky130_fd_sc_hd__o21ai_1
X_12900_ _12928_/A VGND VGND VPWR VPWR _14463_/A sky130_fd_sc_hd__buf_1
XFILLER_47_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12831_ _12831_/A VGND VGND VPWR VPWR _12832_/A sky130_fd_sc_hd__buf_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _15550_/A _15550_/B VGND VGND VPWR VPWR _15690_/B sky130_fd_sc_hd__or2_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12829_/A _12832_/B _10422_/A VGND VGND VPWR VPWR _12762_/Y sky130_fd_sc_hd__o21ai_1
X_15481_ _14790_/A _15452_/B _15452_/X _15480_/X VGND VGND VPWR VPWR _15481_/X sky130_fd_sc_hd__o22a_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14501_/A VGND VGND VPWR VPWR _15211_/A sky130_fd_sc_hd__buf_1
X_11713_ _11713_/A _11720_/B VGND VGND VPWR VPWR _11713_/Y sky130_fd_sc_hd__nor2_1
X_12693_ _10566_/A _12664_/A _10566_/Y _12664_/Y VGND VGND VPWR VPWR _12694_/B sky130_fd_sc_hd__o22a_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _13274_/A _14429_/B _14429_/Y _14431_/X VGND VGND VPWR VPWR _14432_/X sky130_fd_sc_hd__o2bb2a_1
X_11644_ _11643_/Y _11493_/X _11546_/Y VGND VGND VPWR VPWR _11644_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 wbs_dat_i[3] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_4
X_14363_ _11706_/A _14248_/A _14249_/B VGND VGND VPWR VPWR _15774_/A sky130_fd_sc_hd__o21ai_2
X_16102_ _16036_/A _16036_/B _16036_/Y VGND VGND VPWR VPWR _16102_/Y sky130_fd_sc_hd__o21ai_1
Xinput16 wbs_adr_i[8] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_2
X_11575_ _09363_/A _11574_/Y _09365_/X VGND VGND VPWR VPWR _11576_/B sky130_fd_sc_hd__o21a_1
X_14294_ _14309_/A _14294_/B VGND VGND VPWR VPWR _15972_/A sky130_fd_sc_hd__or2_1
X_13314_ _14771_/A _13303_/B _13303_/Y VGND VGND VPWR VPWR _13314_/Y sky130_fd_sc_hd__o21ai_1
X_10526_ _10514_/Y _10524_/X _10525_/Y VGND VGND VPWR VPWR _10526_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16033_ _16022_/Y _16031_/X _16032_/Y VGND VGND VPWR VPWR _16033_/X sky130_fd_sc_hd__o21a_1
X_13245_ _14733_/A _13288_/B VGND VGND VPWR VPWR _13245_/Y sky130_fd_sc_hd__nor2_1
X_10457_ _09122_/A _10456_/X _09122_/A _10456_/X VGND VGND VPWR VPWR _11213_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_124_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13176_ _14564_/A _13103_/B _13103_/Y VGND VGND VPWR VPWR _13176_/Y sky130_fd_sc_hd__o21ai_1
X_10388_ _10451_/A _12698_/A _10387_/Y VGND VGND VPWR VPWR _10388_/X sky130_fd_sc_hd__a21o_1
X_12127_ _12050_/X _12126_/Y _12050_/X _12126_/Y VGND VGND VPWR VPWR _12139_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12058_ _12026_/Y _12056_/X _12057_/Y VGND VGND VPWR VPWR _12058_/X sky130_fd_sc_hd__o21a_1
X_11009_ _12852_/A VGND VGND VPWR VPWR _15063_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15817_ _15817_/A _15817_/B VGND VGND VPWR VPWR _15817_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15748_ _15676_/X _15747_/Y _15676_/X _15747_/Y VGND VGND VPWR VPWR _15809_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15679_ _15679_/A _15679_/B VGND VGND VPWR VPWR _15679_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08984_ _08984_/A _08984_/B VGND VGND VPWR VPWR _11460_/B sky130_fd_sc_hd__or2_1
XFILLER_102_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09605_ _09510_/X _09604_/X _09510_/X _09604_/X VGND VGND VPWR VPWR _09980_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09536_ _09549_/A _09549_/B VGND VGND VPWR VPWR _09613_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09467_ _10014_/A _09467_/B VGND VGND VPWR VPWR _09467_/X sky130_fd_sc_hd__or2_1
XFILLER_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08418_ _08418_/A VGND VGND VPWR VPWR _08418_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09398_ _12854_/A VGND VGND VPWR VPWR _15060_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08349_ _08349_/A VGND VGND VPWR VPWR _08349_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11360_ _12303_/A VGND VGND VPWR VPWR _14132_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10311_ _10309_/A _10309_/B _10310_/A _10309_/Y _10310_/Y VGND VGND VPWR VPWR _10367_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13030_ _14669_/A _13030_/B VGND VGND VPWR VPWR _13030_/X sky130_fd_sc_hd__or2_1
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11291_ _09785_/A _09785_/B _09785_/Y VGND VGND VPWR VPWR _11291_/X sky130_fd_sc_hd__o21a_1
XFILLER_121_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10242_ _10242_/A _10242_/B VGND VGND VPWR VPWR _10242_/X sky130_fd_sc_hd__or2_1
XFILLER_79_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10173_ _10248_/A _10173_/B VGND VGND VPWR VPWR _10173_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14981_ _14980_/Y _14945_/X _14942_/Y VGND VGND VPWR VPWR _14981_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13932_ _15392_/A _13940_/B VGND VGND VPWR VPWR _14041_/A sky130_fd_sc_hd__and2_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13863_ _13777_/X _13794_/A _13793_/X VGND VGND VPWR VPWR _13863_/X sky130_fd_sc_hd__o21a_1
X_15602_ _15602_/A VGND VGND VPWR VPWR _15602_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13794_ _13794_/A _13793_/X VGND VGND VPWR VPWR _13794_/X sky130_fd_sc_hd__or2b_1
X_12814_ _12769_/A _12769_/B _12769_/Y VGND VGND VPWR VPWR _12814_/Y sky130_fd_sc_hd__o21ai_1
X_15533_ _15478_/X _15532_/Y _15478_/X _15532_/Y VGND VGND VPWR VPWR _15616_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12745_ _12696_/A _12696_/B _12696_/Y VGND VGND VPWR VPWR _12745_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15464_ _15464_/A _15464_/B VGND VGND VPWR VPWR _15464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12676_/A VGND VGND VPWR VPWR _12676_/Y sky130_fd_sc_hd__inv_2
X_15395_ _15396_/A _15396_/B VGND VGND VPWR VPWR _15395_/X sky130_fd_sc_hd__or2_1
X_14415_ _11785_/A _14414_/X _11784_/X VGND VGND VPWR VPWR _14416_/A sky130_fd_sc_hd__o21ai_2
X_11627_ _13496_/A _11626_/B _11626_/X _11508_/X VGND VGND VPWR VPWR _11627_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14346_ _13420_/Y _14345_/X _13420_/Y _14345_/X VGND VGND VPWR VPWR _14347_/B sky130_fd_sc_hd__a2bb2oi_1
X_11558_ _13545_/A _11558_/B VGND VGND VPWR VPWR _11558_/X sky130_fd_sc_hd__or2_1
XFILLER_7_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10509_ _09836_/Y _10508_/Y _09836_/A _10508_/A _09941_/A VGND VGND VPWR VPWR _13609_/A
+ sky130_fd_sc_hd__o221a_2
X_16016_ _16036_/A _16036_/B VGND VGND VPWR VPWR _16016_/Y sky130_fd_sc_hd__nor2_1
X_14277_ _14277_/A VGND VGND VPWR VPWR _14277_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11489_ _11587_/A _11489_/B VGND VGND VPWR VPWR _12393_/A sky130_fd_sc_hd__nor2_2
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13228_ _13200_/A _13200_/B _13200_/Y VGND VGND VPWR VPWR _13228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13159_ _13196_/A _13196_/B VGND VGND VPWR VPWR _13159_/Y sky130_fd_sc_hd__nor2_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09321_ _09470_/B _09859_/A _09354_/A VGND VGND VPWR VPWR _09321_/X sky130_fd_sc_hd__o21a_1
X_09252_ _09252_/A _09252_/B VGND VGND VPWR VPWR _10065_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09183_ _09525_/B _09156_/B _09156_/X VGND VGND VPWR VPWR _09184_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08967_ _08682_/X _08966_/X _08682_/X _08966_/X VGND VGND VPWR VPWR _11393_/A sky130_fd_sc_hd__o2bb2a_1
X_08898_ _08685_/X _08897_/X _08685_/X _08897_/X VGND VGND VPWR VPWR _08974_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10860_ _09418_/A _09418_/B _09418_/Y VGND VGND VPWR VPWR _10861_/A sky130_fd_sc_hd__o21ai_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09519_ _09518_/A _09518_/B _09563_/A _09518_/X VGND VGND VPWR VPWR _09519_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10791_ _09908_/A _09908_/B _09911_/A VGND VGND VPWR VPWR _10791_/X sky130_fd_sc_hd__o21ba_1
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _12530_/A _12530_/B VGND VGND VPWR VPWR _12530_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12461_ _12462_/A _12459_/X _12460_/X VGND VGND VPWR VPWR _12461_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11412_ _12235_/A VGND VGND VPWR VPWR _14047_/A sky130_fd_sc_hd__inv_2
X_14200_ _14111_/Y _14199_/X _14111_/Y _14199_/X VGND VGND VPWR VPWR _14201_/B sky130_fd_sc_hd__a2bb2oi_1
X_15180_ _15157_/X _15179_/Y _15157_/X _15179_/Y VGND VGND VPWR VPWR _15181_/B sky130_fd_sc_hd__a2bb2o_1
X_14131_ _14132_/A _14133_/A VGND VGND VPWR VPWR _14131_/Y sky130_fd_sc_hd__nor2_1
X_12392_ _12364_/X _12391_/Y _12364_/X _12391_/Y VGND VGND VPWR VPWR _12458_/B sky130_fd_sc_hd__a2bb2o_1
X_11343_ _11492_/A _11342_/Y _11492_/A _11342_/Y VGND VGND VPWR VPWR _11344_/B sky130_fd_sc_hd__a2bb2o_1
X_14062_ _14062_/A _14062_/B VGND VGND VPWR VPWR _14062_/X sky130_fd_sc_hd__or2_1
X_11274_ _12858_/A VGND VGND VPWR VPWR _15054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13013_ _14497_/A _13013_/B VGND VGND VPWR VPWR _13013_/X sky130_fd_sc_hd__or2_1
X_10225_ _10224_/A _10224_/B _10309_/A VGND VGND VPWR VPWR _10226_/A sky130_fd_sc_hd__o21bai_1
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10156_ _10115_/A _10115_/B _10116_/A VGND VGND VPWR VPWR _10159_/A sky130_fd_sc_hd__a21bo_1
X_14964_ _15563_/A _14982_/B VGND VGND VPWR VPWR _14964_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10087_ _10087_/A _10087_/B VGND VGND VPWR VPWR _11520_/B sky130_fd_sc_hd__or2_1
X_13915_ _14623_/A _13848_/B _13848_/Y VGND VGND VPWR VPWR _13915_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14895_ _15524_/A _14910_/B VGND VGND VPWR VPWR _14895_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13846_ _14627_/A _13846_/B VGND VGND VPWR VPWR _13846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13777_ _13704_/X _13721_/A _13720_/X VGND VGND VPWR VPWR _13777_/X sky130_fd_sc_hd__o21a_1
X_10989_ _10954_/X _10988_/X _10954_/X _10988_/X VGND VGND VPWR VPWR _11128_/B sky130_fd_sc_hd__a2bb2o_1
X_15516_ _15519_/A _15519_/B VGND VGND VPWR VPWR _15639_/A sky130_fd_sc_hd__and2_1
X_12728_ _12718_/X _12727_/X _12718_/X _12727_/X VGND VGND VPWR VPWR _12783_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15447_ _15447_/A _15412_/X VGND VGND VPWR VPWR _15447_/X sky130_fd_sc_hd__or2b_1
X_12659_ _10369_/Y _12658_/Y _10307_/Y VGND VGND VPWR VPWR _12660_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15378_ _15378_/A _15339_/X VGND VGND VPWR VPWR _15378_/X sky130_fd_sc_hd__or2b_1
XFILLER_129_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14329_ _14335_/A _14329_/B VGND VGND VPWR VPWR _15958_/A sky130_fd_sc_hd__or2_1
X_09870_ _09450_/Y _09869_/X _09474_/X VGND VGND VPWR VPWR _09870_/X sky130_fd_sc_hd__o21a_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08821_ _09221_/A _09456_/B _08716_/X VGND VGND VPWR VPWR _08822_/A sky130_fd_sc_hd__o21ai_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _10008_/A _10134_/A VGND VGND VPWR VPWR _08752_/X sky130_fd_sc_hd__or2_1
XFILLER_66_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08683_ _09547_/A _08622_/A _08624_/Y _08682_/X VGND VGND VPWR VPWR _08683_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09304_ _09304_/A _10235_/A VGND VGND VPWR VPWR _09304_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09235_ _09235_/A _09681_/A VGND VGND VPWR VPWR _09629_/A sky130_fd_sc_hd__or2_1
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09166_ _10009_/B _09166_/B VGND VGND VPWR VPWR _09167_/B sky130_fd_sc_hd__or2_1
XFILLER_119_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09097_ _09070_/A _09070_/B _09071_/B VGND VGND VPWR VPWR _09409_/A sky130_fd_sc_hd__a21bo_1
XFILLER_89_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10010_ _10010_/A _10010_/B VGND VGND VPWR VPWR _10038_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09999_ _09999_/A _09999_/B VGND VGND VPWR VPWR _10000_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11961_ _11959_/X _11960_/Y _11959_/X _11960_/Y VGND VGND VPWR VPWR _11962_/B sky130_fd_sc_hd__a2bb2o_1
X_10912_ _14631_/A _10883_/B _10883_/X _10911_/X VGND VGND VPWR VPWR _10912_/X sky130_fd_sc_hd__o22a_1
X_13700_ _13730_/A _13698_/X _13699_/X VGND VGND VPWR VPWR _13700_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14680_ _15184_/A _14681_/B VGND VGND VPWR VPWR _14682_/A sky130_fd_sc_hd__and2_1
X_11892_ _11892_/A _11892_/B VGND VGND VPWR VPWR _11892_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10843_ _13058_/A _10842_/B _10842_/Y VGND VGND VPWR VPWR _10843_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13631_ _13596_/Y _13628_/Y _13630_/Y VGND VGND VPWR VPWR _13632_/A sky130_fd_sc_hd__o21ai_1
X_16350_ _08230_/X _16468_/Q _08233_/X _16349_/X _16343_/X VGND VGND VPWR VPWR _16468_/D
+ sky130_fd_sc_hd__o221a_2
X_10774_ _13073_/A _10720_/B _10720_/Y _10773_/X VGND VGND VPWR VPWR _10774_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13562_ _15032_/A _13525_/B _13525_/Y VGND VGND VPWR VPWR _13562_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16281_ _16338_/A _16338_/B VGND VGND VPWR VPWR _16281_/Y sky130_fd_sc_hd__nor2_1
X_12513_ _13444_/A _11363_/B _11363_/Y VGND VGND VPWR VPWR _12514_/B sky130_fd_sc_hd__o21a_1
X_15301_ _15280_/X _15300_/Y _15280_/X _15300_/Y VGND VGND VPWR VPWR _15347_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13493_ _11618_/Y _12379_/A _11535_/Y _13492_/X VGND VGND VPWR VPWR _13493_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15232_ _15178_/A _15178_/B _15178_/Y VGND VGND VPWR VPWR _15232_/Y sky130_fd_sc_hd__o21ai_1
X_12444_ _12444_/A VGND VGND VPWR VPWR _13973_/A sky130_fd_sc_hd__buf_1
XFILLER_8_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15163_ _15163_/A _15163_/B VGND VGND VPWR VPWR _15163_/Y sky130_fd_sc_hd__nor2_1
X_12375_ _11319_/A _12270_/A _11518_/B VGND VGND VPWR VPWR _12375_/Y sky130_fd_sc_hd__a21oi_1
X_14114_ _14114_/A VGND VGND VPWR VPWR _14880_/A sky130_fd_sc_hd__inv_2
X_15094_ _15069_/A _15069_/B _15069_/Y _15093_/X VGND VGND VPWR VPWR _15094_/X sky130_fd_sc_hd__a2bb2o_1
X_11326_ _11326_/A VGND VGND VPWR VPWR _11326_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14045_ _14430_/A _13938_/B _14430_/A _13938_/B VGND VGND VPWR VPWR _14045_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11257_ _11449_/A _11212_/B _11212_/Y _11256_/X VGND VGND VPWR VPWR _11257_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11188_ _14060_/A _11188_/B VGND VGND VPWR VPWR _11188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10208_ _10287_/A VGND VGND VPWR VPWR _10903_/A sky130_fd_sc_hd__inv_2
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10139_ _10139_/A _10139_/B VGND VGND VPWR VPWR _10139_/Y sky130_fd_sc_hd__nor2_1
X_15996_ _15970_/A _15970_/B _15970_/Y VGND VGND VPWR VPWR _15996_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14947_ _14948_/A _14948_/B VGND VGND VPWR VPWR _14949_/A sky130_fd_sc_hd__and2_1
XFILLER_63_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14878_ _14823_/X _14877_/X _14823_/X _14877_/X VGND VGND VPWR VPWR _14920_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13829_ _13829_/A VGND VGND VPWR VPWR _14646_/A sky130_fd_sc_hd__inv_2
XFILLER_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09020_ _09470_/A _08567_/X _09020_/S VGND VGND VPWR VPWR _09555_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09922_ _09923_/A _09923_/B VGND VGND VPWR VPWR _11298_/B sky130_fd_sc_hd__and2_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09853_ _09853_/A _09853_/B VGND VGND VPWR VPWR _09897_/A sky130_fd_sc_hd__and2_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08804_ _09250_/A VGND VGND VPWR VPWR _09494_/A sky130_fd_sc_hd__buf_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _09785_/A _09785_/B VGND VGND VPWR VPWR _09784_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08735_ _08712_/Y _08733_/Y _08734_/X VGND VGND VPWR VPWR _08736_/A sky130_fd_sc_hd__o21ai_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _08934_/A _09232_/B _09232_/A _08398_/Y VGND VGND VPWR VPWR _08667_/A sky130_fd_sc_hd__o22a_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08597_ _08597_/A _10114_/B VGND VGND VPWR VPWR _08598_/A sky130_fd_sc_hd__or2_1
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10490_ _10490_/A VGND VGND VPWR VPWR _10490_/Y sky130_fd_sc_hd__inv_2
X_09218_ _09803_/A VGND VGND VPWR VPWR _09696_/A sky130_fd_sc_hd__inv_2
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09149_ _09518_/A _09148_/X _08521_/B VGND VGND VPWR VPWR _09150_/S sky130_fd_sc_hd__o21ba_1
XFILLER_107_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12160_ _12160_/A _12160_/B VGND VGND VPWR VPWR _12160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11111_ _09993_/A _09662_/B _09662_/Y VGND VGND VPWR VPWR _11111_/X sky130_fd_sc_hd__o21a_1
X_12091_ _12779_/A _12168_/A _12090_/Y VGND VGND VPWR VPWR _12091_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11042_ _12842_/A VGND VGND VPWR VPWR _15078_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15850_ _14178_/A _15849_/X _12635_/X VGND VGND VPWR VPWR _15850_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14801_ _14728_/X _14800_/X _14728_/X _14800_/X VGND VGND VPWR VPWR _14802_/B sky130_fd_sc_hd__a2bb2o_1
X_15781_ _15781_/A _15781_/B VGND VGND VPWR VPWR _16241_/A sky130_fd_sc_hd__or2_1
X_12993_ _13015_/A _13016_/B VGND VGND VPWR VPWR _13085_/A sky130_fd_sc_hd__and2_1
XFILLER_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14732_ _14796_/A _14730_/X _14731_/X VGND VGND VPWR VPWR _14732_/X sky130_fd_sc_hd__o21a_1
X_11944_ _11903_/A _11943_/Y _11903_/A _11943_/Y VGND VGND VPWR VPWR _11972_/B sky130_fd_sc_hd__a2bb2o_1
X_14663_ _14610_/Y _14661_/X _14662_/Y VGND VGND VPWR VPWR _14663_/X sky130_fd_sc_hd__o21a_1
X_11875_ _11840_/X _11874_/Y _11840_/X _11874_/Y VGND VGND VPWR VPWR _11901_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16402_ _16402_/A _16402_/B VGND VGND VPWR VPWR _16402_/X sky130_fd_sc_hd__or2_1
X_13614_ _12914_/A _14430_/B _12914_/A _14430_/B VGND VGND VPWR VPWR _13614_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10826_ _10826_/A _10826_/B VGND VGND VPWR VPWR _10826_/Y sky130_fd_sc_hd__nand2_1
X_14594_ _14529_/A _14529_/B _14526_/X _14529_/Y VGND VGND VPWR VPWR _14594_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16333_ _16290_/Y _16331_/X _16332_/Y VGND VGND VPWR VPWR _16333_/X sky130_fd_sc_hd__o21a_1
X_13545_ _13545_/A VGND VGND VPWR VPWR _15420_/A sky130_fd_sc_hd__buf_1
X_10757_ _13753_/A VGND VGND VPWR VPWR _11958_/A sky130_fd_sc_hd__inv_2
X_16264_ _16264_/A _16264_/B VGND VGND VPWR VPWR _16264_/Y sky130_fd_sc_hd__nand2_1
X_13476_ _13450_/A _13450_/B _13450_/Y VGND VGND VPWR VPWR _13476_/X sky130_fd_sc_hd__o21a_1
X_10688_ _10688_/A _10688_/B VGND VGND VPWR VPWR _10688_/Y sky130_fd_sc_hd__nand2_1
X_15215_ _15216_/A _15216_/B VGND VGND VPWR VPWR _15268_/A sky130_fd_sc_hd__and2_1
X_12427_ _12424_/X _12426_/X _12424_/X _12426_/X VGND VGND VPWR VPWR _12429_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16195_ _16106_/A _15807_/B _15807_/Y VGND VGND VPWR VPWR _16196_/A sky130_fd_sc_hd__o21ai_1
XFILLER_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12358_ _13204_/A _12358_/B VGND VGND VPWR VPWR _12358_/Y sky130_fd_sc_hd__nor2_1
X_15146_ _15146_/A _15146_/B VGND VGND VPWR VPWR _15146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12289_ _12253_/X _12288_/Y _12253_/X _12288_/Y VGND VGND VPWR VPWR _12358_/B sky130_fd_sc_hd__a2bb2o_1
X_15077_ _15031_/X _15076_/X _15031_/X _15076_/X VGND VGND VPWR VPWR _15078_/B sky130_fd_sc_hd__a2bb2o_1
X_11309_ _11312_/A VGND VGND VPWR VPWR _11309_/Y sky130_fd_sc_hd__inv_2
X_14028_ _14028_/A _14028_/B VGND VGND VPWR VPWR _14028_/X sky130_fd_sc_hd__and2_1
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15979_ _15909_/Y _15978_/Y _15912_/Y VGND VGND VPWR VPWR _15979_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08520_ _09476_/B VGND VGND VPWR VPWR _08694_/A sky130_fd_sc_hd__buf_1
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08451_ _08710_/A VGND VGND VPWR VPWR _09332_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08382_ _08366_/A _08365_/Y _08366_/Y _08365_/A _08419_/A VGND VGND VPWR VPWR _08642_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09003_ _11569_/A _09003_/B VGND VGND VPWR VPWR _12300_/A sky130_fd_sc_hd__or2_1
XFILLER_129_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09905_ _09857_/A _09857_/B _09904_/Y VGND VGND VPWR VPWR _10653_/A sky130_fd_sc_hd__a21oi_1
XFILLER_100_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _09836_/A VGND VGND VPWR VPWR _09836_/Y sky130_fd_sc_hd__inv_2
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09767_ _09730_/A _09730_/B _09733_/A VGND VGND VPWR VPWR _10052_/A sky130_fd_sc_hd__a21bo_1
XFILLER_27_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08718_ _08718_/A _09462_/B VGND VGND VPWR VPWR _08718_/Y sky130_fd_sc_hd__nor2_1
X_09698_ _09698_/A _09698_/B VGND VGND VPWR VPWR _09730_/A sky130_fd_sc_hd__or2_1
XFILLER_27_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08649_ input2/X input18/X _08392_/Y _08481_/Y _08392_/A VGND VGND VPWR VPWR _08650_/B
+ sky130_fd_sc_hd__o32a_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11559_/A _11472_/X _11558_/X VGND VGND VPWR VPWR _11685_/A sky130_fd_sc_hd__o21ai_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10611_ _10524_/X _10610_/Y _10524_/X _10610_/Y VGND VGND VPWR VPWR _10629_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11591_ _09864_/X _09933_/X _09864_/X _09933_/X VGND VGND VPWR VPWR _11592_/B sky130_fd_sc_hd__a2bb2oi_1
X_13330_ _13287_/A _13329_/Y _13287_/A _13329_/Y VGND VGND VPWR VPWR _13331_/B sky130_fd_sc_hd__a2bb2o_1
X_10542_ _10541_/A _10541_/B _10541_/Y _09393_/A VGND VGND VPWR VPWR _11021_/A sky130_fd_sc_hd__o211a_1
X_13261_ _13926_/A VGND VGND VPWR VPWR _14725_/A sky130_fd_sc_hd__inv_2
XFILLER_6_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12212_ _14021_/A _12212_/B VGND VGND VPWR VPWR _12212_/Y sky130_fd_sc_hd__nand2_1
X_15000_ _11751_/A _14999_/X _11750_/X VGND VGND VPWR VPWR _15000_/X sky130_fd_sc_hd__o21a_1
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10473_ _10469_/Y _10471_/A _10469_/A _10471_/Y _10982_/A VGND VGND VPWR VPWR _11852_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13192_ _13192_/A _13192_/B VGND VGND VPWR VPWR _13192_/Y sky130_fd_sc_hd__nand2_1
X_12143_ _13918_/A _12143_/B VGND VGND VPWR VPWR _12143_/X sky130_fd_sc_hd__or2_1
X_12074_ _13584_/A _12073_/B _12073_/X _11984_/X VGND VGND VPWR VPWR _12074_/X sky130_fd_sc_hd__o22a_1
X_15902_ _15902_/A _15902_/B VGND VGND VPWR VPWR _15902_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11025_ _11025_/A _10916_/X VGND VGND VPWR VPWR _11025_/X sky130_fd_sc_hd__or2b_1
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15833_ _16192_/A VGND VGND VPWR VPWR _16160_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15764_ _14907_/X _15763_/X _14907_/X _15763_/X VGND VGND VPWR VPWR _15765_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14715_ _15392_/A VGND VGND VPWR VPWR _15398_/A sky130_fd_sc_hd__buf_1
X_12976_ _12935_/X _12975_/Y _12935_/X _12975_/Y VGND VGND VPWR VPWR _13024_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15695_ _15689_/Y _15693_/Y _15694_/Y VGND VGND VPWR VPWR _15695_/X sky130_fd_sc_hd__o21a_1
X_11927_ _11990_/B _11926_/X _11990_/B _11926_/X VGND VGND VPWR VPWR _11986_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14646_ _14646_/A _14646_/B VGND VGND VPWR VPWR _14646_/X sky130_fd_sc_hd__or2_1
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11858_ _11859_/A _11859_/B VGND VGND VPWR VPWR _11860_/A sky130_fd_sc_hd__and2_1
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14577_ _14563_/Y _14575_/X _14576_/Y VGND VGND VPWR VPWR _14577_/X sky130_fd_sc_hd__o21a_1
X_11789_ _12829_/A _11717_/B _11717_/Y VGND VGND VPWR VPWR _11789_/Y sky130_fd_sc_hd__a21oi_1
X_10809_ _10809_/A _11925_/A VGND VGND VPWR VPWR _10809_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16316_ _16316_/A _16316_/B VGND VGND VPWR VPWR _16316_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13528_ _13528_/A _13528_/B VGND VGND VPWR VPWR _13528_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16247_ _16241_/A _16246_/A _16241_/Y _16246_/Y _16247_/C1 VGND VGND VPWR VPWR _16248_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13459_ _13458_/Y _12786_/X _12722_/Y VGND VGND VPWR VPWR _13459_/X sky130_fd_sc_hd__o21a_1
X_16178_ _16264_/A _16330_/A VGND VGND VPWR VPWR _16178_/Y sky130_fd_sc_hd__nor2_1
X_15129_ _15072_/A _15072_/B _15072_/Y VGND VGND VPWR VPWR _15129_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09621_ _09972_/A VGND VGND VPWR VPWR _09960_/A sky130_fd_sc_hd__buf_1
XFILLER_28_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09552_ _09607_/A _09550_/X _09607_/B VGND VGND VPWR VPWR _09552_/X sky130_fd_sc_hd__o21ba_1
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08503_ _08701_/A _08503_/B VGND VGND VPWR VPWR _09448_/B sky130_fd_sc_hd__or2_2
X_09483_ _08765_/A _09475_/X _08765_/A _09475_/X VGND VGND VPWR VPWR _09484_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08434_ _08434_/A VGND VGND VPWR VPWR _08434_/Y sky130_fd_sc_hd__inv_2
X_08365_ _08365_/A VGND VGND VPWR VPWR _08365_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08296_ _08296_/A VGND VGND VPWR VPWR _08296_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09819_ _09819_/A _09819_/B VGND VGND VPWR VPWR _09820_/B sky130_fd_sc_hd__or2_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12830_ _12829_/A _12829_/B _12829_/Y VGND VGND VPWR VPWR _12830_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12761_ _10342_/X _10424_/B _10342_/X _10424_/B VGND VGND VPWR VPWR _12832_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15480_ _14794_/A _15455_/B _15455_/X _15479_/Y VGND VGND VPWR VPWR _15480_/X sky130_fd_sc_hd__o22a_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _15208_/A _14512_/B VGND VGND VPWR VPWR _14561_/A sky130_fd_sc_hd__and2_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12692_/A _12692_/B VGND VGND VPWR VPWR _12692_/Y sky130_fd_sc_hd__nor2_1
X_11712_ _10210_/A _10347_/A _10284_/Y _13479_/B _11721_/B VGND VGND VPWR VPWR _11720_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _15396_/A _14430_/B _10428_/X _14430_/X VGND VGND VPWR VPWR _14431_/X sky130_fd_sc_hd__o22a_1
X_11643_ _12390_/A _11643_/B VGND VGND VPWR VPWR _11643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput28 wbs_dat_i[4] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__buf_4
XFILLER_128_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16101_ _16101_/A _16104_/B VGND VGND VPWR VPWR _16101_/Y sky130_fd_sc_hd__nor2_1
X_14362_ _14368_/A _14362_/B VGND VGND VPWR VPWR _14364_/A sky130_fd_sc_hd__nor2_1
Xinput17 wbs_adr_i[9] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_1
X_11574_ _11574_/A VGND VGND VPWR VPWR _11574_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14293_ _13447_/X _14292_/X _13447_/X _14292_/X VGND VGND VPWR VPWR _14294_/B sky130_fd_sc_hd__a2bb2oi_1
X_13313_ _13313_/A _13313_/B VGND VGND VPWR VPWR _13313_/X sky130_fd_sc_hd__and2_1
X_10525_ _11835_/A _10525_/B VGND VGND VPWR VPWR _10525_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16032_ _16032_/A _16032_/B VGND VGND VPWR VPWR _16032_/Y sky130_fd_sc_hd__nand2_1
X_13244_ _13193_/X _13243_/Y _13193_/X _13243_/Y VGND VGND VPWR VPWR _13288_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10456_ _09418_/A _09123_/B _09123_/Y VGND VGND VPWR VPWR _10456_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13175_ _13829_/A VGND VGND VPWR VPWR _15331_/A sky130_fd_sc_hd__buf_1
XFILLER_6_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12126_ _12037_/A _12051_/B _12051_/Y VGND VGND VPWR VPWR _12126_/Y sky130_fd_sc_hd__o21ai_1
X_10387_ _10451_/A _11803_/A VGND VGND VPWR VPWR _10387_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12057_ _12057_/A _12057_/B VGND VGND VPWR VPWR _12057_/Y sky130_fd_sc_hd__nand2_1
X_11008_ _13584_/A VGND VGND VPWR VPWR _12852_/A sky130_fd_sc_hd__buf_1
XFILLER_38_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15816_ _15731_/Y _15814_/X _15815_/Y VGND VGND VPWR VPWR _15816_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15747_ _15677_/A _15677_/B _15677_/Y VGND VGND VPWR VPWR _15747_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12959_ _14757_/A _12944_/B _12944_/Y VGND VGND VPWR VPWR _12959_/Y sky130_fd_sc_hd__o21ai_1
X_15678_ _15614_/Y _15676_/X _15677_/Y VGND VGND VPWR VPWR _15678_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14629_ _14579_/X _14628_/Y _14579_/X _14628_/Y VGND VGND VPWR VPWR _14652_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08983_ _08880_/X _08981_/X _09001_/B VGND VGND VPWR VPWR _08983_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ _09494_/A _09494_/B _09494_/Y VGND VGND VPWR VPWR _09604_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09535_ _09551_/A _09551_/B VGND VGND VPWR VPWR _09607_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09466_ _10015_/A _08597_/A _09455_/Y _09465_/X VGND VGND VPWR VPWR _09466_/X sky130_fd_sc_hd__o22a_1
X_08417_ _08351_/Y _08413_/Y _10016_/A VGND VGND VPWR VPWR _08417_/Y sky130_fd_sc_hd__a21oi_1
X_09397_ _13649_/A VGND VGND VPWR VPWR _12854_/A sky130_fd_sc_hd__buf_1
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08348_ _08348_/A VGND VGND VPWR VPWR _08348_/Y sky130_fd_sc_hd__inv_2
X_08279_ input9/X _08279_/B VGND VGND VPWR VPWR _08279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11290_ _11288_/Y _11289_/Y _11167_/Y VGND VGND VPWR VPWR _11492_/A sky130_fd_sc_hd__o21ai_1
X_10310_ _10310_/A VGND VGND VPWR VPWR _10310_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10241_ _10241_/A _10241_/B VGND VGND VPWR VPWR _10241_/X sky130_fd_sc_hd__or2_1
XFILLER_121_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10172_ _10124_/A _10124_/B _10125_/B VGND VGND VPWR VPWR _10173_/B sky130_fd_sc_hd__a21bo_1
XFILLER_78_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14980_ _15425_/A _14980_/B VGND VGND VPWR VPWR _14980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13931_ _13839_/X _13930_/Y _13839_/X _13930_/Y VGND VGND VPWR VPWR _13940_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13862_ _13776_/X _13798_/A _13797_/X VGND VGND VPWR VPWR _13862_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15601_ _15601_/A VGND VGND VPWR VPWR _15601_/Y sky130_fd_sc_hd__inv_2
X_13793_ _13793_/A _13793_/B VGND VGND VPWR VPWR _13793_/X sky130_fd_sc_hd__or2_1
X_12813_ _12846_/A _12846_/B VGND VGND VPWR VPWR _12813_/Y sky130_fd_sc_hd__nor2_1
X_15532_ _15458_/A _15458_/B _15458_/Y VGND VGND VPWR VPWR _15532_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12773_/A _12773_/B VGND VGND VPWR VPWR _12744_/Y sky130_fd_sc_hd__nor2_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15463_ _15401_/X _15462_/X _15401_/X _15462_/X VGND VGND VPWR VPWR _15464_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _11518_/Y _12674_/Y _11324_/Y VGND VGND VPWR VPWR _12676_/A sky130_fd_sc_hd__o21ai_2
X_15394_ _12043_/A _15393_/Y _12043_/A _15393_/Y VGND VGND VPWR VPWR _15396_/B sky130_fd_sc_hd__a2bb2o_1
X_14414_ _12832_/A _11717_/B _14413_/X VGND VGND VPWR VPWR _14414_/X sky130_fd_sc_hd__o21a_1
X_11626_ _11626_/A _11626_/B VGND VGND VPWR VPWR _11626_/X sky130_fd_sc_hd__and2_1
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14345_ _14096_/A _13421_/B _13421_/Y VGND VGND VPWR VPWR _14345_/X sky130_fd_sc_hd__o21a_1
X_11557_ _13545_/A _11558_/B VGND VGND VPWR VPWR _11559_/A sky130_fd_sc_hd__and2_1
XFILLER_116_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10508_ _10508_/A VGND VGND VPWR VPWR _10508_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16015_ _15953_/X _16014_/X _15953_/X _16014_/X VGND VGND VPWR VPWR _16036_/B sky130_fd_sc_hd__a2bb2o_1
X_14276_ _14186_/Y _14274_/Y _14275_/Y VGND VGND VPWR VPWR _14277_/A sky130_fd_sc_hd__o21ai_1
X_11488_ _09665_/X _11487_/X _09665_/X _11487_/X VGND VGND VPWR VPWR _11489_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13227_ _14597_/A VGND VGND VPWR VPWR _14739_/A sky130_fd_sc_hd__buf_1
X_10439_ _10439_/A VGND VGND VPWR VPWR _10439_/Y sky130_fd_sc_hd__inv_2
X_13158_ _13114_/X _13157_/Y _13114_/X _13157_/Y VGND VGND VPWR VPWR _13196_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13089_ _13747_/A VGND VGND VPWR VPWR _15264_/A sky130_fd_sc_hd__buf_1
X_12109_ _12062_/X _12108_/Y _12062_/X _12108_/Y VGND VGND VPWR VPWR _12151_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09320_ _09531_/A _09737_/A VGND VGND VPWR VPWR _09354_/A sky130_fd_sc_hd__or2_1
XFILLER_34_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09251_ _09456_/A _09251_/B VGND VGND VPWR VPWR _10069_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09182_ _09430_/A _09185_/B VGND VGND VPWR VPWR _09182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08966_ _09547_/A _08622_/A _08624_/A VGND VGND VPWR VPWR _08966_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08897_ _09553_/A _08584_/A _08586_/A VGND VGND VPWR VPWR _08897_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09518_ _09518_/A _09518_/B VGND VGND VPWR VPWR _09518_/X sky130_fd_sc_hd__and2_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10790_ _10789_/Y _10652_/X _10698_/Y VGND VGND VPWR VPWR _10790_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09449_ _09482_/A _09525_/A VGND VGND VPWR VPWR _09449_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12460_ _15285_/A _12460_/B VGND VGND VPWR VPWR _12460_/X sky130_fd_sc_hd__or2_1
XFILLER_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11411_ _11411_/A _11411_/B _12232_/B VGND VGND VPWR VPWR _12235_/A sky130_fd_sc_hd__or3_1
X_12391_ _12953_/A _12454_/B _12390_/Y VGND VGND VPWR VPWR _12391_/Y sky130_fd_sc_hd__o21ai_1
X_14130_ _14061_/X _14129_/X _14061_/X _14129_/X VGND VGND VPWR VPWR _14133_/A sky130_fd_sc_hd__a2bb2o_1
X_11342_ _13793_/A _11491_/B _11341_/Y VGND VGND VPWR VPWR _11342_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14061_ _14123_/A _14059_/X _14060_/X VGND VGND VPWR VPWR _14061_/X sky130_fd_sc_hd__o21a_1
X_11273_ _11273_/A VGND VGND VPWR VPWR _12858_/A sky130_fd_sc_hd__buf_1
XFILLER_4_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13012_ _13012_/A VGND VGND VPWR VPWR _14497_/A sky130_fd_sc_hd__buf_1
X_10224_ _10224_/A _10224_/B VGND VGND VPWR VPWR _10309_/A sky130_fd_sc_hd__and2_1
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10155_ _10155_/A _10155_/B VGND VGND VPWR VPWR _10155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14963_ _14933_/Y _14962_/Y _14933_/Y _14962_/Y VGND VGND VPWR VPWR _14982_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10086_ _10040_/X _10084_/X _11316_/B VGND VGND VPWR VPWR _10086_/X sky130_fd_sc_hd__o21a_1
X_14894_ _14818_/X _14893_/X _14818_/X _14893_/X VGND VGND VPWR VPWR _14910_/B sky130_fd_sc_hd__a2bb2o_1
X_13914_ _13914_/A VGND VGND VPWR VPWR _15406_/A sky130_fd_sc_hd__buf_1
XFILLER_90_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13845_ _13824_/Y _13843_/X _13844_/Y VGND VGND VPWR VPWR _13845_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13776_ _13801_/A _13774_/X _13775_/X VGND VGND VPWR VPWR _13776_/X sky130_fd_sc_hd__o21a_1
X_10988_ _13507_/A _11130_/B _13507_/A _11130_/B VGND VGND VPWR VPWR _10988_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15515_ _15512_/A _15512_/B _15512_/X _15651_/A VGND VGND VPWR VPWR _15519_/B sky130_fd_sc_hd__o22a_1
X_12727_ _12684_/A _12684_/B _12684_/Y VGND VGND VPWR VPWR _12727_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15446_ _15446_/A _15446_/B VGND VGND VPWR VPWR _15446_/X sky130_fd_sc_hd__and2_1
XFILLER_90_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12658_ _10224_/A _10224_/B _12657_/Y VGND VGND VPWR VPWR _12658_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11609_ _11609_/A _12423_/B VGND VGND VPWR VPWR _11609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12589_ _12589_/A VGND VGND VPWR VPWR _12589_/Y sky130_fd_sc_hd__inv_2
X_15377_ _15408_/A _15408_/B VGND VGND VPWR VPWR _15453_/A sky130_fd_sc_hd__and2_1
X_14328_ _13435_/Y _14327_/X _13435_/Y _14327_/X VGND VGND VPWR VPWR _14329_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_7_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14259_ _14259_/A VGND VGND VPWR VPWR _14259_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08820_ _09252_/A VGND VGND VPWR VPWR _09498_/A sky130_fd_sc_hd__buf_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _09339_/B VGND VGND VPWR VPWR _10134_/A sky130_fd_sc_hd__buf_1
X_08682_ _09538_/A _08635_/A _08637_/Y _08681_/Y VGND VGND VPWR VPWR _08682_/X sky130_fd_sc_hd__o22a_1
XFILLER_66_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09303_ _09304_/A _10235_/A VGND VGND VPWR VPWR _09303_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09234_ _09707_/B VGND VGND VPWR VPWR _09681_/A sky130_fd_sc_hd__inv_2
XFILLER_22_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09165_ _10010_/B _09165_/B VGND VGND VPWR VPWR _09166_/B sky130_fd_sc_hd__or2_1
XFILLER_107_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09096_ _09716_/A VGND VGND VPWR VPWR _09717_/A sky130_fd_sc_hd__buf_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09998_ _09964_/X _11510_/A _11509_/B VGND VGND VPWR VPWR _09999_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08949_ _09459_/B VGND VGND VPWR VPWR _09539_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11960_ _13001_/A _11890_/B _11890_/Y VGND VGND VPWR VPWR _11960_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10911_ _13825_/A _10891_/B _10891_/Y _10910_/X VGND VGND VPWR VPWR _10911_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11891_ _11959_/A _11889_/Y _11890_/Y VGND VGND VPWR VPWR _11891_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10842_ _12066_/A _10842_/B VGND VGND VPWR VPWR _10842_/Y sky130_fd_sc_hd__nand2_1
X_13630_ _15131_/A _13630_/B VGND VGND VPWR VPWR _13630_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10773_ _13078_/A _10729_/B _10729_/Y _10772_/X VGND VGND VPWR VPWR _10773_/X sky130_fd_sc_hd__a2bb2o_1
X_13561_ _13561_/A VGND VGND VPWR VPWR _13561_/Y sky130_fd_sc_hd__inv_2
X_16280_ _16271_/X _16279_/Y _16271_/X _16279_/Y VGND VGND VPWR VPWR _16338_/B sky130_fd_sc_hd__o2bb2a_1
X_12512_ _14132_/A VGND VGND VPWR VPWR _13444_/A sky130_fd_sc_hd__buf_1
X_15300_ _14665_/A _15243_/B _15243_/Y VGND VGND VPWR VPWR _15300_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15231_ _15285_/A _15285_/B VGND VGND VPWR VPWR _15287_/A sky130_fd_sc_hd__nor2_1
X_13492_ _11513_/Y _12273_/A _11331_/Y _13491_/X VGND VGND VPWR VPWR _13492_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12443_ _12443_/A VGND VGND VPWR VPWR _15285_/A sky130_fd_sc_hd__buf_1
XFILLER_60_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15162_ _12419_/A _15161_/Y _12419_/A _15161_/Y VGND VGND VPWR VPWR _15163_/B sky130_fd_sc_hd__a2bb2o_1
X_12374_ _12684_/A _12373_/B _12373_/X _12273_/B VGND VGND VPWR VPWR _12417_/B sky130_fd_sc_hd__a22o_1
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14113_ _14108_/Y _14111_/Y _14112_/Y VGND VGND VPWR VPWR _14113_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15093_ _15072_/A _15072_/B _15072_/Y _15092_/X VGND VGND VPWR VPWR _15093_/X sky130_fd_sc_hd__a2bb2o_1
X_11325_ _11518_/A _11518_/B _11324_/Y VGND VGND VPWR VPWR _11326_/A sky130_fd_sc_hd__o21ai_2
XFILLER_109_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14044_ _14048_/A VGND VGND VPWR VPWR _14815_/A sky130_fd_sc_hd__buf_1
X_11256_ _14028_/A _11218_/B _11218_/Y _11255_/X VGND VGND VPWR VPWR _11256_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11187_ _11092_/X _11186_/X _11092_/X _11186_/X VGND VGND VPWR VPWR _11188_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10207_ _10346_/B VGND VGND VPWR VPWR _10463_/A sky130_fd_sc_hd__clkbuf_2
X_15995_ _16055_/A _16055_/B VGND VGND VPWR VPWR _16059_/A sky130_fd_sc_hd__and2_1
XFILLER_94_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10138_ _10133_/A _10133_/B _10134_/B VGND VGND VPWR VPWR _10139_/B sky130_fd_sc_hd__a21bo_1
XFILLER_94_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14946_ _14943_/Y _14945_/X _14943_/Y _14945_/X VGND VGND VPWR VPWR _14948_/B sky130_fd_sc_hd__a2bb2o_1
X_10069_ _10069_/A _10069_/B VGND VGND VPWR VPWR _10069_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14877_ _14786_/A _14786_/B _14786_/A _14786_/B VGND VGND VPWR VPWR _14877_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13828_ _14635_/A _13842_/B VGND VGND VPWR VPWR _13828_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13759_ _15264_/A _13759_/B VGND VGND VPWR VPWR _13759_/X sky130_fd_sc_hd__or2_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15429_ _15424_/Y _15428_/X _15424_/Y _15428_/X VGND VGND VPWR VPWR _15429_/X sky130_fd_sc_hd__a2bb2o_1
X_09921_ _09921_/A _09920_/Y VGND VGND VPWR VPWR _09923_/B sky130_fd_sc_hd__or2b_1
XFILLER_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09852_ _09853_/A _09853_/B VGND VGND VPWR VPWR _09855_/A sky130_fd_sc_hd__nor2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08803_ _10014_/A _09249_/B VGND VGND VPWR VPWR _08803_/Y sky130_fd_sc_hd__nor2_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _10083_/A _09781_/Y _09782_/Y VGND VGND VPWR VPWR _09785_/B sky130_fd_sc_hd__o21ai_1
XFILLER_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08734_ _10012_/A _09531_/A VGND VGND VPWR VPWR _08734_/X sky130_fd_sc_hd__or2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _08665_/A VGND VGND VPWR VPWR _08671_/A sky130_fd_sc_hd__inv_2
XFILLER_26_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08596_ _08596_/A VGND VGND VPWR VPWR _10114_/B sky130_fd_sc_hd__inv_2
XFILLER_26_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09217_ _09217_/A _09217_/B VGND VGND VPWR VPWR _09803_/A sky130_fd_sc_hd__or2_2
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09148_ _08762_/A _09147_/X _08532_/B VGND VGND VPWR VPWR _09148_/X sky130_fd_sc_hd__o21ba_1
X_09079_ _10011_/B _09078_/B _09165_/B VGND VGND VPWR VPWR _09760_/A sky130_fd_sc_hd__a21bo_1
X_11110_ _13053_/A _10998_/B _10998_/Y _10929_/X VGND VGND VPWR VPWR _11110_/X sky130_fd_sc_hd__a2bb2o_1
X_12090_ _12779_/A _12168_/A VGND VGND VPWR VPWR _12090_/Y sky130_fd_sc_hd__nor2_1
X_11041_ _13564_/A VGND VGND VPWR VPWR _12842_/A sky130_fd_sc_hd__buf_1
XFILLER_1_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14800_ _14800_/A _14729_/X VGND VGND VPWR VPWR _14800_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15780_ _15774_/A _16028_/A _15656_/A _16028_/B VGND VGND VPWR VPWR _15781_/B sky130_fd_sc_hd__a22o_1
XFILLER_76_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12992_ _12927_/X _12991_/Y _12927_/X _12991_/Y VGND VGND VPWR VPWR _13016_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14731_ _14731_/A _14731_/B VGND VGND VPWR VPWR _14731_/X sky130_fd_sc_hd__or2_1
X_11943_ _13695_/A _11904_/B _11904_/Y VGND VGND VPWR VPWR _11943_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14662_ _15347_/A _14662_/B VGND VGND VPWR VPWR _14662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11874_ _13625_/A _11841_/B _11841_/Y VGND VGND VPWR VPWR _11874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16401_ _16394_/Y _16398_/Y _16399_/Y _16400_/Y VGND VGND VPWR VPWR _16401_/X sky130_fd_sc_hd__o211a_1
X_13613_ _10421_/B _11789_/Y _10424_/B _11791_/B VGND VGND VPWR VPWR _14430_/B sky130_fd_sc_hd__o22a_1
XFILLER_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10825_ _09263_/B _10242_/B _10242_/X VGND VGND VPWR VPWR _10826_/B sky130_fd_sc_hd__a21boi_1
X_16332_ _16332_/A _16332_/B VGND VGND VPWR VPWR _16332_/Y sky130_fd_sc_hd__nand2_1
X_14593_ _14532_/A _14532_/B _14525_/X _14532_/Y VGND VGND VPWR VPWR _14593_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10756_ _10761_/A _10756_/B VGND VGND VPWR VPWR _13753_/A sky130_fd_sc_hd__or2_1
X_13544_ _13458_/A _13495_/B _13495_/X _13543_/X VGND VGND VPWR VPWR _13544_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16263_ _16186_/Y _16261_/X _16262_/Y VGND VGND VPWR VPWR _16263_/X sky130_fd_sc_hd__o21a_1
X_13475_ _14335_/A VGND VGND VPWR VPWR _14309_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10687_ _09269_/B _10243_/B _10243_/X VGND VGND VPWR VPWR _10688_/B sky130_fd_sc_hd__a21boi_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16194_ _16260_/A _16326_/A VGND VGND VPWR VPWR _16194_/Y sky130_fd_sc_hd__nor2_1
X_15214_ _10522_/Y _15213_/Y _10522_/Y _15213_/Y VGND VGND VPWR VPWR _15216_/B sky130_fd_sc_hd__o2bb2a_1
X_12426_ _12426_/A _12426_/B VGND VGND VPWR VPWR _12426_/X sky130_fd_sc_hd__or2_1
X_15145_ _12835_/X _15144_/X _12835_/X _15144_/X VGND VGND VPWR VPWR _15146_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12357_ _12295_/A _12248_/X _12294_/X VGND VGND VPWR VPWR _12357_/X sky130_fd_sc_hd__o21a_1
X_12288_ _13042_/A _12360_/B _12287_/Y VGND VGND VPWR VPWR _12288_/Y sky130_fd_sc_hd__o21ai_1
X_15076_ _15076_/A _15032_/X VGND VGND VPWR VPWR _15076_/X sky130_fd_sc_hd__or2b_1
X_11308_ _11307_/A _11307_/B _11307_/Y _10957_/X VGND VGND VPWR VPWR _11506_/A sky130_fd_sc_hd__o211a_1
X_11239_ _12230_/A VGND VGND VPWR VPWR _13349_/A sky130_fd_sc_hd__buf_1
X_14027_ _13947_/X _14026_/Y _13947_/X _14026_/Y VGND VGND VPWR VPWR _14028_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15978_ _15978_/A _15978_/B VGND VGND VPWR VPWR _15978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14929_ _14863_/Y _14927_/X _14928_/Y VGND VGND VPWR VPWR _14929_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08450_ _10010_/A VGND VGND VPWR VPWR _08710_/A sky130_fd_sc_hd__inv_2
X_08381_ _08401_/A VGND VGND VPWR VPWR _08419_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09002_ _08981_/X _09001_/X _08981_/X _09001_/X VGND VGND VPWR VPWR _09003_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09904_ _09904_/A VGND VGND VPWR VPWR _09904_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _09799_/A _09799_/B _09834_/Y VGND VGND VPWR VPWR _09836_/A sky130_fd_sc_hd__a21oi_1
XFILLER_112_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09766_ _09766_/A VGND VGND VPWR VPWR _09776_/A sky130_fd_sc_hd__inv_2
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08717_ _08717_/A _08717_/B VGND VGND VPWR VPWR _08717_/X sky130_fd_sc_hd__or2_1
X_09697_ _08592_/A _09728_/B _08592_/A _09728_/B VGND VGND VPWR VPWR _09698_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08648_ _09230_/A _10110_/B VGND VGND VPWR VPWR _08648_/X sky130_fd_sc_hd__or2_1
XFILLER_27_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08579_ _09209_/B VGND VGND VPWR VPWR _08579_/Y sky130_fd_sc_hd__inv_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10610_ _11835_/A _10525_/B _10525_/Y VGND VGND VPWR VPWR _10610_/Y sky130_fd_sc_hd__o21ai_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11590_ _11590_/A _11590_/B VGND VGND VPWR VPWR _12452_/A sky130_fd_sc_hd__or2_2
X_10541_ _10541_/A _10541_/B VGND VGND VPWR VPWR _10541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13260_ _14727_/A _13279_/B VGND VGND VPWR VPWR _13260_/Y sky130_fd_sc_hd__nor2_1
X_12211_ _12148_/X _12210_/X _12148_/X _12210_/X VGND VGND VPWR VPWR _12212_/B sky130_fd_sc_hd__a2bb2o_1
X_10472_ _10472_/A VGND VGND VPWR VPWR _10982_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13191_ _13168_/Y _13189_/X _13190_/Y VGND VGND VPWR VPWR _13191_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12142_ _12222_/A _12140_/X _12141_/X VGND VGND VPWR VPWR _12142_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12073_ _13584_/A _12073_/B VGND VGND VPWR VPWR _12073_/X sky130_fd_sc_hd__and2_1
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15901_ _15862_/Y _15899_/X _15900_/Y VGND VGND VPWR VPWR _15901_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11024_ _15069_/A VGND VGND VPWR VPWR _13910_/A sky130_fd_sc_hd__buf_1
XFILLER_77_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15832_ _15832_/A VGND VGND VPWR VPWR _16192_/A sky130_fd_sc_hd__buf_1
XFILLER_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15763_ _14908_/A _14908_/B _14908_/Y VGND VGND VPWR VPWR _15763_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12975_ _14477_/A _12936_/B _12936_/Y VGND VGND VPWR VPWR _12975_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14714_ _14725_/A _14725_/B VGND VGND VPWR VPWR _14807_/A sky130_fd_sc_hd__nor2_1
X_11926_ _11926_/A _11925_/X VGND VGND VPWR VPWR _11926_/X sky130_fd_sc_hd__or2b_1
X_15694_ _15694_/A _15694_/B VGND VGND VPWR VPWR _15694_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14645_ _14644_/A _14644_/B _11065_/B _14644_/Y VGND VGND VPWR VPWR _14645_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11857_ _10566_/A _11856_/A _10566_/Y _11920_/B VGND VGND VPWR VPWR _11859_/B sky130_fd_sc_hd__o22a_1
X_14576_ _14576_/A _14576_/B VGND VGND VPWR VPWR _14576_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11788_ _11788_/A VGND VGND VPWR VPWR _12829_/A sky130_fd_sc_hd__buf_1
X_10808_ _11990_/A VGND VGND VPWR VPWR _11925_/A sky130_fd_sc_hd__inv_2
X_16315_ _16316_/A _16316_/B VGND VGND VPWR VPWR _16315_/Y sky130_fd_sc_hd__nor2_1
X_13527_ _10326_/X _13482_/X _10326_/X _13482_/X VGND VGND VPWR VPWR _13528_/B sky130_fd_sc_hd__o2bb2a_1
X_10739_ _09958_/A _09640_/B _09640_/Y VGND VGND VPWR VPWR _10741_/A sky130_fd_sc_hd__o21ai_1
X_16246_ _16246_/A VGND VGND VPWR VPWR _16246_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13458_ _13458_/A _13458_/B VGND VGND VPWR VPWR _13458_/Y sky130_fd_sc_hd__nor2_1
X_16177_ _16264_/B VGND VGND VPWR VPWR _16330_/A sky130_fd_sc_hd__buf_1
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12409_ _12409_/A _12409_/B VGND VGND VPWR VPWR _12409_/Y sky130_fd_sc_hd__nand2_1
X_13389_ _13364_/X _13388_/X _13364_/X _13388_/X VGND VGND VPWR VPWR _13440_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15128_ _15128_/A _15128_/B VGND VGND VPWR VPWR _15128_/Y sky130_fd_sc_hd__nand2_1
X_15059_ _15043_/X _15058_/X _15043_/X _15058_/X VGND VGND VPWR VPWR _15060_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09620_ _09507_/X _09619_/X _09507_/X _09619_/X VGND VGND VPWR VPWR _09972_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09551_ _09551_/A _09551_/B VGND VGND VPWR VPWR _09607_/B sky130_fd_sc_hd__and2_1
XFILLER_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08502_ _08308_/Y _08501_/A _08308_/A _08501_/Y VGND VGND VPWR VPWR _08503_/B sky130_fd_sc_hd__o22a_1
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09482_ _09482_/A _09482_/B VGND VGND VPWR VPWR _09482_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08433_ _09209_/B _08428_/X _09324_/A VGND VGND VPWR VPWR _08433_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08364_ _08364_/A _08364_/B VGND VGND VPWR VPWR _08365_/A sky130_fd_sc_hd__or2_1
X_08295_ input22/X _08306_/B _08307_/A _08309_/A VGND VGND VPWR VPWR _08296_/A sky130_fd_sc_hd__o22a_1
XFILLER_117_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09818_ _09818_/A _09818_/B VGND VGND VPWR VPWR _09819_/B sky130_fd_sc_hd__or2_1
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09749_ _10034_/A VGND VGND VPWR VPWR _09749_/X sky130_fd_sc_hd__buf_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12760_ _12763_/A _12763_/B VGND VGND VPWR VPWR _12760_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12691_ _10685_/A _12666_/A _10685_/Y _12666_/Y VGND VGND VPWR VPWR _12692_/B sky130_fd_sc_hd__o22a_1
X_11711_ _11711_/A _11711_/B VGND VGND VPWR VPWR _11721_/B sky130_fd_sc_hd__or2_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A _14430_/B VGND VGND VPWR VPWR _14430_/X sky130_fd_sc_hd__and2_1
X_11642_ _12452_/A _11641_/B _11641_/X VGND VGND VPWR VPWR _11642_/X sky130_fd_sc_hd__a21bo_1
XFILLER_42_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14361_ _14378_/A _14378_/B VGND VGND VPWR VPWR _14361_/Y sky130_fd_sc_hd__nor2_1
X_16100_ _16096_/Y _16098_/X _16099_/Y VGND VGND VPWR VPWR _16104_/B sky130_fd_sc_hd__o21ai_1
X_11573_ _15437_/A _11561_/B _11561_/Y _11466_/X VGND VGND VPWR VPWR _11573_/Y sky130_fd_sc_hd__a2bb2oi_1
X_13312_ _13305_/A _13311_/Y _13305_/A _13311_/Y VGND VGND VPWR VPWR _13313_/B sky130_fd_sc_hd__a2bb2o_1
Xinput18 wbs_dat_i[0] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_2
Xinput29 wbs_dat_i[5] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_4
X_14292_ _13448_/A _13448_/B _13448_/Y VGND VGND VPWR VPWR _14292_/X sky130_fd_sc_hd__o21a_1
X_10524_ _13610_/A _10523_/B _10522_/Y _10523_/Y VGND VGND VPWR VPWR _10524_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16031_ _16025_/Y _16029_/X _16030_/Y VGND VGND VPWR VPWR _16031_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13243_ _13194_/A _13194_/B _13194_/Y VGND VGND VPWR VPWR _13243_/Y sky130_fd_sc_hd__o21ai_1
X_10455_ _10455_/A VGND VGND VPWR VPWR _10966_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13174_ _13825_/A _13186_/B VGND VGND VPWR VPWR _13174_/Y sky130_fd_sc_hd__nor2_1
X_12125_ _13922_/A _12141_/B VGND VGND VPWR VPWR _12222_/A sky130_fd_sc_hd__and2_1
XFILLER_69_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10386_ _11803_/A VGND VGND VPWR VPWR _12698_/A sky130_fd_sc_hd__buf_1
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12056_ _12030_/Y _12054_/X _12055_/Y VGND VGND VPWR VPWR _12056_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11007_ _11007_/A VGND VGND VPWR VPWR _13584_/A sky130_fd_sc_hd__buf_1
X_15815_ _16114_/A _15815_/B VGND VGND VPWR VPWR _15815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15746_ _15752_/A _15746_/B VGND VGND VPWR VPWR _16108_/A sky130_fd_sc_hd__nor2_1
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12958_ _13793_/A VGND VGND VPWR VPWR _14749_/A sky130_fd_sc_hd__inv_2
XFILLER_46_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15677_ _15677_/A _15677_/B VGND VGND VPWR VPWR _15677_/Y sky130_fd_sc_hd__nand2_1
X_11909_ _13633_/A _11909_/B VGND VGND VPWR VPWR _11909_/Y sky130_fd_sc_hd__nor2_1
X_12889_ _12848_/A _12848_/B _12848_/Y VGND VGND VPWR VPWR _12889_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14628_ _14580_/A _14580_/B _14580_/Y VGND VGND VPWR VPWR _14628_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14559_ _14578_/A _14578_/B VGND VGND VPWR VPWR _14559_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16229_ _16227_/A _16228_/A _16227_/Y _16228_/Y _15832_/A VGND VGND VPWR VPWR _16251_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08982_ _08982_/A _08982_/B VGND VGND VPWR VPWR _09001_/B sky130_fd_sc_hd__or2_1
XFILLER_130_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09603_ _09984_/A _09656_/B VGND VGND VPWR VPWR _09603_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09534_ _09553_/A _09553_/B VGND VGND VPWR VPWR _09601_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09465_ _10016_/A _08610_/A _09456_/Y _09464_/X VGND VGND VPWR VPWR _09465_/X sky130_fd_sc_hd__o22a_1
X_08416_ _09221_/A VGND VGND VPWR VPWR _10016_/A sky130_fd_sc_hd__buf_1
XFILLER_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09396_ _09396_/A VGND VGND VPWR VPWR _13649_/A sky130_fd_sc_hd__buf_1
X_08347_ _08347_/A _08347_/B VGND VGND VPWR VPWR _08348_/A sky130_fd_sc_hd__or2_1
X_08278_ _08278_/A VGND VGND VPWR VPWR _08279_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10240_ _10240_/A _10240_/B VGND VGND VPWR VPWR _10240_/X sky130_fd_sc_hd__or2_1
XFILLER_106_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10171_ _10111_/A _10111_/B _10112_/A VGND VGND VPWR VPWR _10248_/A sky130_fd_sc_hd__a21bo_1
XFILLER_120_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13930_ _14646_/A _13840_/B _13840_/Y VGND VGND VPWR VPWR _13930_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15600_ _15600_/A _15542_/X VGND VGND VPWR VPWR _15601_/A sky130_fd_sc_hd__or2b_1
X_13861_ _13800_/Y _13859_/X _13860_/Y VGND VGND VPWR VPWR _13861_/X sky130_fd_sc_hd__o21a_1
X_13792_ _13793_/A _13793_/B VGND VGND VPWR VPWR _13794_/A sky130_fd_sc_hd__and2_1
XFILLER_62_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12812_ _12770_/X _12811_/Y _12770_/X _12811_/Y VGND VGND VPWR VPWR _12846_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15531_ _15534_/A _15534_/B VGND VGND VPWR VPWR _15531_/Y sky130_fd_sc_hd__nor2_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12713_/X _12742_/X _12713_/X _12742_/X VGND VGND VPWR VPWR _12773_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15462_ _15462_/A _15402_/X VGND VGND VPWR VPWR _15462_/X sky130_fd_sc_hd__or2b_1
XFILLER_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _10424_/A _10421_/B _12832_/A _11717_/B VGND VGND VPWR VPWR _14413_/X sky130_fd_sc_hd__a22o_1
X_12674_ _12674_/A VGND VGND VPWR VPWR _12674_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15393_ _15329_/A _15329_/B _15329_/Y VGND VGND VPWR VPWR _15393_/Y sky130_fd_sc_hd__a21oi_1
X_11625_ _12410_/A _11624_/B _11624_/Y VGND VGND VPWR VPWR _11625_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14344_ _14256_/A _14343_/Y _14256_/A _14343_/Y VGND VGND VPWR VPWR _14382_/A sky130_fd_sc_hd__a2bb2o_1
X_11556_ _11481_/X _11555_/X _11481_/X _11555_/X VGND VGND VPWR VPWR _11558_/B sky130_fd_sc_hd__a2bb2o_1
X_14275_ _15857_/A _14275_/B VGND VGND VPWR VPWR _14275_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10507_ _09832_/A _09832_/B _09833_/A VGND VGND VPWR VPWR _10508_/A sky130_fd_sc_hd__o21ai_1
X_16014_ _16014_/A _15954_/X VGND VGND VPWR VPWR _16014_/X sky130_fd_sc_hd__or2b_1
X_13226_ _15060_/A VGND VGND VPWR VPWR _14597_/A sky130_fd_sc_hd__inv_2
X_11487_ _09997_/A _09666_/B _09666_/Y VGND VGND VPWR VPWR _11487_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10438_ _10438_/A VGND VGND VPWR VPWR _10438_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13157_ _15249_/A _13115_/B _13115_/Y VGND VGND VPWR VPWR _13157_/Y sky130_fd_sc_hd__o21ai_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _11759_/A _10369_/B VGND VGND VPWR VPWR _10369_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13088_ _13088_/A VGND VGND VPWR VPWR _13747_/A sky130_fd_sc_hd__inv_2
X_12108_ _13198_/A _12063_/B _12063_/Y VGND VGND VPWR VPWR _12108_/Y sky130_fd_sc_hd__o21ai_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12039_ _11963_/X _12038_/X _11963_/X _12038_/X VGND VGND VPWR VPWR _12049_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15729_ _15683_/A _15683_/B _15683_/Y VGND VGND VPWR VPWR _15729_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09250_ _09250_/A _10127_/A VGND VGND VPWR VPWR _10073_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09181_ _09177_/Y _09179_/Y _09180_/Y VGND VGND VPWR VPWR _09185_/B sky130_fd_sc_hd__o21ai_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08965_ _08968_/A _08968_/B VGND VGND VPWR VPWR _08965_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08896_ _08976_/A _08976_/B VGND VGND VPWR VPWR _08896_/X sky130_fd_sc_hd__and2_1
XFILLER_84_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09517_ _09482_/A _09482_/B _09482_/Y _09516_/X VGND VGND VPWR VPWR _09563_/A sky130_fd_sc_hd__o2bb2a_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09448_ _09448_/A _09448_/B VGND VGND VPWR VPWR _09448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09379_ _09355_/X _09378_/X _09355_/X _09378_/X VGND VGND VPWR VPWR _09380_/A sky130_fd_sc_hd__a2bb2o_1
X_11410_ _12320_/A VGND VGND VPWR VPWR _13406_/A sky130_fd_sc_hd__inv_2
X_12390_ _12390_/A _12454_/B VGND VGND VPWR VPWR _12390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11341_ _12362_/A _11491_/B VGND VGND VPWR VPWR _11341_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14060_ _14060_/A _14060_/B VGND VGND VPWR VPWR _14060_/X sky130_fd_sc_hd__or2_1
X_11272_ _13786_/A VGND VGND VPWR VPWR _11273_/A sky130_fd_sc_hd__buf_1
XFILLER_121_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13011_ _13000_/Y _13009_/X _13010_/Y VGND VGND VPWR VPWR _13011_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10223_ _10175_/Y _10222_/A _10175_/A _10222_/Y _10463_/A VGND VGND VPWR VPWR _10224_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10154_ _08793_/B _10129_/B _10130_/B VGND VGND VPWR VPWR _10155_/B sky130_fd_sc_hd__a21bo_1
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14962_ _14971_/A _14971_/B _14961_/Y VGND VGND VPWR VPWR _14962_/Y sky130_fd_sc_hd__o21ai_1
X_10085_ _10085_/A _10085_/B VGND VGND VPWR VPWR _11316_/B sky130_fd_sc_hd__or2_1
X_14893_ _14806_/A _14806_/B _14806_/A _14806_/B VGND VGND VPWR VPWR _14893_/X sky130_fd_sc_hd__a2bb2o_1
X_13913_ _15408_/A _13950_/B VGND VGND VPWR VPWR _13913_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13844_ _14631_/A _13844_/B VGND VGND VPWR VPWR _13844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13775_ _13775_/A _13775_/B VGND VGND VPWR VPWR _13775_/X sky130_fd_sc_hd__or2_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10987_ _10963_/X _10986_/X _10963_/X _10986_/X VGND VGND VPWR VPWR _11130_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15514_ _15474_/X _15513_/Y _15474_/X _15513_/Y VGND VGND VPWR VPWR _15651_/A sky130_fd_sc_hd__a2bb2o_1
X_12726_ _12785_/A _12785_/B VGND VGND VPWR VPWR _12726_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15445_ _15413_/X _15444_/X _15413_/X _15444_/X VGND VGND VPWR VPWR _15446_/B sky130_fd_sc_hd__a2bb2o_1
X_12657_ _10201_/Y _12656_/Y _10213_/Y VGND VGND VPWR VPWR _12657_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15376_ _15340_/X _15375_/X _15340_/X _15375_/X VGND VGND VPWR VPWR _15408_/B sky130_fd_sc_hd__a2bb2o_1
X_11608_ _10122_/Y _11607_/A _10237_/B _11607_/Y _11526_/A VGND VGND VPWR VPWR _12423_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_129_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ _12585_/Y _12587_/Y _12585_/A _12587_/A _11706_/A VGND VGND VPWR VPWR _12619_/A
+ sky130_fd_sc_hd__o221a_1
X_14327_ _14112_/A _13436_/B _13436_/Y VGND VGND VPWR VPWR _14327_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11539_ _11508_/X _11538_/X _11508_/X _11538_/X VGND VGND VPWR VPWR _11631_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14258_ _14222_/Y _14256_/Y _14257_/Y VGND VGND VPWR VPWR _14259_/A sky130_fd_sc_hd__o21ai_1
XFILLER_131_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14189_ _14207_/A _14189_/B VGND VGND VPWR VPWR _15860_/A sky130_fd_sc_hd__or2_1
X_13209_ _14934_/A _13452_/B VGND VGND VPWR VPWR _13209_/Y sky130_fd_sc_hd__nand2_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08749_/A _08748_/Y _08749_/Y _09341_/B VGND VGND VPWR VPWR _09339_/B sky130_fd_sc_hd__o22a_1
XFILLER_38_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08681_ _09230_/A _10110_/B _08648_/X _08680_/X VGND VGND VPWR VPWR _08681_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_26_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09302_ _09301_/A _08946_/Y _09301_/Y _08946_/A VGND VGND VPWR VPWR _10235_/A sky130_fd_sc_hd__o22a_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09233_ _09678_/A VGND VGND VPWR VPWR _09707_/B sky130_fd_sc_hd__clkbuf_2
X_09164_ _08765_/Y _09158_/A _08765_/A _09158_/Y VGND VGND VPWR VPWR _10010_/B sky130_fd_sc_hd__o22a_1
XFILLER_21_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09095_ _10018_/B _09071_/B _09072_/B VGND VGND VPWR VPWR _09716_/A sky130_fd_sc_hd__a21bo_1
XFILLER_103_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09997_ _09997_/A _09997_/B VGND VGND VPWR VPWR _11509_/B sky130_fd_sc_hd__or2_1
XFILLER_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08948_ _08952_/A _08952_/B VGND VGND VPWR VPWR _08948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08879_ _08878_/Y _08866_/X _08878_/Y _08866_/X VGND VGND VPWR VPWR _08982_/B sky130_fd_sc_hd__o2bb2a_1
X_10910_ _10898_/Y _10908_/X _10909_/Y VGND VGND VPWR VPWR _10910_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11890_ _13001_/A _11890_/B VGND VGND VPWR VPWR _11890_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10841_ _10936_/A _10840_/Y _10936_/A _10840_/Y VGND VGND VPWR VPWR _10842_/B sky130_fd_sc_hd__a2bb2o_1
X_10772_ _13083_/A _10738_/B _10738_/Y _10771_/X VGND VGND VPWR VPWR _10772_/X sky130_fd_sc_hd__a2bb2o_1
X_13560_ _13560_/A _13560_/B VGND VGND VPWR VPWR _13561_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12511_ _12637_/A _12637_/B VGND VGND VPWR VPWR _14284_/A sky130_fd_sc_hd__and2_1
X_13491_ _11309_/Y _12179_/A _11157_/Y _13490_/X VGND VGND VPWR VPWR _13491_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15230_ _15175_/Y _15229_/Y _15175_/Y _15229_/Y VGND VGND VPWR VPWR _15285_/B sky130_fd_sc_hd__a2bb2o_1
X_12442_ _13463_/A _12439_/B _12439_/X _12441_/X VGND VGND VPWR VPWR _12442_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15161_ _15161_/A VGND VGND VPWR VPWR _15161_/Y sky130_fd_sc_hd__inv_2
X_12373_ _12373_/A _12373_/B VGND VGND VPWR VPWR _12373_/X sky130_fd_sc_hd__or2_1
XFILLER_126_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14112_ _14112_/A _14112_/B VGND VGND VPWR VPWR _14112_/Y sky130_fd_sc_hd__nand2_1
X_15092_ _15075_/A _15075_/B _15075_/Y _15091_/X VGND VGND VPWR VPWR _15092_/X sky130_fd_sc_hd__a2bb2o_1
X_11324_ _11518_/A _11518_/B VGND VGND VPWR VPWR _11324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14043_ _14043_/A _14043_/B VGND VGND VPWR VPWR _14043_/Y sky130_fd_sc_hd__nor2_1
X_11255_ _14032_/A _11224_/B _11224_/Y _11254_/X VGND VGND VPWR VPWR _11255_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10206_ _10206_/A VGND VGND VPWR VPWR _11721_/A sky130_fd_sc_hd__inv_2
XFILLER_121_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11186_ _11186_/A _11093_/X VGND VGND VPWR VPWR _11186_/X sky130_fd_sc_hd__or2b_1
XFILLER_79_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15994_ _15971_/X _15993_/X _15971_/X _15993_/X VGND VGND VPWR VPWR _16055_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10137_ _10139_/A VGND VGND VPWR VPWR _10238_/B sky130_fd_sc_hd__buf_1
X_14945_ _14837_/X _14944_/Y _14844_/Y VGND VGND VPWR VPWR _14945_/X sky130_fd_sc_hd__o21a_1
X_10068_ _10067_/A _10067_/B _09971_/A _10067_/X VGND VGND VPWR VPWR _10071_/A sky130_fd_sc_hd__a22o_1
XFILLER_63_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14876_ _14876_/A VGND VGND VPWR VPWR _15544_/A sky130_fd_sc_hd__buf_1
XFILLER_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13827_ _13758_/X _13826_/X _13758_/X _13826_/X VGND VGND VPWR VPWR _13842_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13758_ _13750_/Y _13756_/X _13757_/Y VGND VGND VPWR VPWR _13758_/X sky130_fd_sc_hd__o21a_1
X_12709_ _12706_/A _12706_/B _12706_/Y _12708_/X VGND VGND VPWR VPWR _12709_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13689_ _14497_/A _13689_/B VGND VGND VPWR VPWR _13689_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15428_ _15426_/X _15427_/Y _15426_/X _15427_/Y VGND VGND VPWR VPWR _15428_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15359_ _15420_/A _15420_/B VGND VGND VPWR VPWR _15435_/A sky130_fd_sc_hd__and2_1
XFILLER_116_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09920_ _09918_/A _09918_/B _09919_/Y VGND VGND VPWR VPWR _09920_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09851_ _09851_/A _09850_/Y VGND VGND VPWR VPWR _09853_/B sky130_fd_sc_hd__or2b_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08802_ _10128_/A VGND VGND VPWR VPWR _09249_/B sky130_fd_sc_hd__buf_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09782_/A _09782_/B VGND VGND VPWR VPWR _09782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08733_ _08733_/A VGND VGND VPWR VPWR _08733_/Y sky130_fd_sc_hd__inv_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08664_ _08665_/A VGND VGND VPWR VPWR _08664_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08595_ _08715_/B VGND VGND VPWR VPWR _08597_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09216_ _09216_/A VGND VGND VPWR VPWR _09216_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09147_ _08770_/A _09015_/X _08543_/B VGND VGND VPWR VPWR _09147_/X sky130_fd_sc_hd__o21ba_1
X_09078_ _10011_/B _09078_/B VGND VGND VPWR VPWR _09165_/B sky130_fd_sc_hd__or2_1
XFILLER_123_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11040_ _13918_/A _11083_/B VGND VGND VPWR VPWR _11222_/A sky130_fd_sc_hd__and2_1
XFILLER_89_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12991_ _14463_/A _12928_/B _12928_/Y VGND VGND VPWR VPWR _12991_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14730_ _14800_/A _14728_/X _14729_/X VGND VGND VPWR VPWR _14730_/X sky130_fd_sc_hd__o21a_1
X_11942_ _11942_/A _11974_/B VGND VGND VPWR VPWR _11942_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14661_ _14614_/Y _14659_/X _14660_/Y VGND VGND VPWR VPWR _14661_/X sky130_fd_sc_hd__o21a_1
X_11873_ _11904_/A _11904_/B VGND VGND VPWR VPWR _11873_/Y sky130_fd_sc_hd__nor2_1
X_16400_ _16407_/D VGND VGND VPWR VPWR _16400_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14592_ _14592_/A VGND VGND VPWR VPWR _15187_/A sky130_fd_sc_hd__buf_1
X_13612_ _13612_/A VGND VGND VPWR VPWR _13612_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10824_ _10812_/X _10823_/Y _10812_/X _10823_/Y VGND VGND VPWR VPWR _10962_/A sky130_fd_sc_hd__o2bb2a_1
X_16331_ _16293_/Y _16329_/X _16330_/Y VGND VGND VPWR VPWR _16331_/X sky130_fd_sc_hd__o21a_1
X_13543_ _15104_/A _13498_/B _13498_/Y _13542_/X VGND VGND VPWR VPWR _13543_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10755_ _11964_/A _10769_/B VGND VGND VPWR VPWR _10896_/A sky130_fd_sc_hd__and2_1
XFILLER_40_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16262_ _16262_/A _16262_/B VGND VGND VPWR VPWR _16262_/Y sky130_fd_sc_hd__nand2_1
X_13474_ _14353_/A VGND VGND VPWR VPWR _14335_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10686_ _10674_/X _10685_/Y _10674_/X _10685_/Y VGND VGND VPWR VPWR _10809_/A sky130_fd_sc_hd__o2bb2a_1
X_16193_ _16260_/B VGND VGND VPWR VPWR _16326_/A sky130_fd_sc_hd__buf_1
X_15213_ _15146_/A _15146_/B _15146_/Y VGND VGND VPWR VPWR _15213_/Y sky130_fd_sc_hd__o21ai_1
X_12425_ _12425_/A VGND VGND VPWR VPWR _12426_/A sky130_fd_sc_hd__inv_2
X_12356_ _14064_/A _12297_/B _12297_/Y _12247_/X VGND VGND VPWR VPWR _12356_/X sky130_fd_sc_hd__a2bb2o_1
X_15144_ _15144_/A _15087_/X VGND VGND VPWR VPWR _15144_/X sky130_fd_sc_hd__or2b_1
XFILLER_114_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11307_ _11307_/A _11307_/B VGND VGND VPWR VPWR _11307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12287_ _12360_/A _12360_/B VGND VGND VPWR VPWR _12287_/Y sky130_fd_sc_hd__nand2_1
X_15075_ _15075_/A _15075_/B VGND VGND VPWR VPWR _15075_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11238_ _14043_/A VGND VGND VPWR VPWR _12230_/A sky130_fd_sc_hd__inv_2
X_14026_ _15406_/A _13948_/B _13948_/Y VGND VGND VPWR VPWR _14026_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11169_ _11289_/A _11168_/Y _11289_/A _11168_/Y VGND VGND VPWR VPWR _11170_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15977_ _15984_/A _15984_/B _15976_/Y VGND VGND VPWR VPWR _15977_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14928_ _15552_/A _14928_/B VGND VGND VPWR VPWR _14928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14859_ _14859_/A _14858_/X VGND VGND VPWR VPWR _14859_/X sky130_fd_sc_hd__or2b_1
XFILLER_63_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08380_ _08662_/A VGND VGND VPWR VPWR _08401_/A sky130_fd_sc_hd__inv_2
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09001_ _08880_/X _09001_/B VGND VGND VPWR VPWR _09001_/X sky130_fd_sc_hd__and2b_1
XFILLER_117_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09903_ _09903_/A _09903_/B VGND VGND VPWR VPWR _10654_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09834_ _09834_/A VGND VGND VPWR VPWR _09834_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09765_ _10049_/A VGND VGND VPWR VPWR _10079_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer30 _16240_/B VGND VGND VPWR VPWR _16313_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_73_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08716_ _08716_/A _08716_/B VGND VGND VPWR VPWR _08716_/X sky130_fd_sc_hd__or2_1
X_09696_ _09696_/A _09696_/B VGND VGND VPWR VPWR _09728_/B sky130_fd_sc_hd__or2_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08647_ _08647_/A VGND VGND VPWR VPWR _10110_/B sky130_fd_sc_hd__inv_2
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08578_ _09209_/A VGND VGND VPWR VPWR _10013_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10540_ _09275_/A _09275_/B _09275_/X VGND VGND VPWR VPWR _10541_/B sky130_fd_sc_hd__a21boi_1
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10471_ _10471_/A VGND VGND VPWR VPWR _10471_/Y sky130_fd_sc_hd__inv_2
X_12210_ _12210_/A _12149_/X VGND VGND VPWR VPWR _12210_/X sky130_fd_sc_hd__or2b_1
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13190_ _13190_/A _13190_/B VGND VGND VPWR VPWR _13190_/Y sky130_fd_sc_hd__nand2_1
X_12141_ _13922_/A _12141_/B VGND VGND VPWR VPWR _12141_/X sky130_fd_sc_hd__or2_1
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12072_ _12071_/Y _11982_/X _12005_/Y VGND VGND VPWR VPWR _12072_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15900_ _15900_/A _15900_/B VGND VGND VPWR VPWR _15900_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11023_ _12848_/A VGND VGND VPWR VPWR _15069_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15831_ _16238_/A VGND VGND VPWR VPWR _15832_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15762_ _15765_/A _15762_/B VGND VGND VPWR VPWR _15799_/A sky130_fd_sc_hd__or2_1
X_12974_ _13699_/A VGND VGND VPWR VPWR _14412_/A sky130_fd_sc_hd__inv_2
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14713_ _14647_/Y _14712_/Y _14647_/Y _14712_/Y VGND VGND VPWR VPWR _14725_/B sky130_fd_sc_hd__a2bb2o_1
X_11925_ _11925_/A _11925_/B VGND VGND VPWR VPWR _11925_/X sky130_fd_sc_hd__or2_1
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15693_ _16053_/A VGND VGND VPWR VPWR _15693_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14644_ _14644_/A _14644_/B VGND VGND VPWR VPWR _14644_/Y sky130_fd_sc_hd__nor2_1
X_11856_ _11856_/A VGND VGND VPWR VPWR _11920_/B sky130_fd_sc_hd__inv_2
X_14575_ _14567_/Y _14573_/X _14574_/Y VGND VGND VPWR VPWR _14575_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11787_ _11787_/A _11787_/B VGND VGND VPWR VPWR _11787_/Y sky130_fd_sc_hd__nor2_1
X_10807_ _10809_/A VGND VGND VPWR VPWR _10807_/Y sky130_fd_sc_hd__inv_2
X_16314_ _16248_/Y _16313_/Y _16248_/Y _16313_/Y VGND VGND VPWR VPWR _16316_/B sky130_fd_sc_hd__o2bb2a_1
X_10738_ _11968_/A _10738_/B VGND VGND VPWR VPWR _10738_/Y sky130_fd_sc_hd__nand2_1
X_13526_ _13528_/A VGND VGND VPWR VPWR _15030_/A sky130_fd_sc_hd__buf_1
XFILLER_41_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16245_ _16245_/A _15782_/X VGND VGND VPWR VPWR _16246_/A sky130_fd_sc_hd__or2b_1
X_13457_ _13130_/X _13456_/X _13130_/X _13456_/X VGND VGND VPWR VPWR _13457_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12408_ _13448_/A _12407_/B _12407_/Y VGND VGND VPWR VPWR _12409_/B sky130_fd_sc_hd__o21a_1
X_10669_ _10671_/A VGND VGND VPWR VPWR _10669_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16176_ _16192_/A _16176_/B VGND VGND VPWR VPWR _16264_/B sky130_fd_sc_hd__or2_1
XFILLER_114_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13388_ _13388_/A _13365_/X VGND VGND VPWR VPWR _13388_/X sky130_fd_sc_hd__or2b_1
XFILLER_126_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12339_ _13396_/A _12339_/B VGND VGND VPWR VPWR _12339_/Y sky130_fd_sc_hd__nand2_1
X_15127_ _15093_/X _15126_/Y _15093_/X _15126_/Y VGND VGND VPWR VPWR _15128_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15058_ _15058_/A _15044_/X VGND VGND VPWR VPWR _15058_/X sky130_fd_sc_hd__or2b_1
XFILLER_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14009_ _14009_/A _14064_/B VGND VGND VPWR VPWR _14135_/A sky130_fd_sc_hd__and2_1
XFILLER_95_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09550_ _09613_/A _09548_/X _09613_/B VGND VGND VPWR VPWR _09550_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08501_ _08501_/A VGND VGND VPWR VPWR _08501_/Y sky130_fd_sc_hd__inv_2
X_09481_ _08757_/A _09477_/X _08757_/A _09477_/X VGND VGND VPWR VPWR _09482_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08432_ _08713_/A VGND VGND VPWR VPWR _09324_/A sky130_fd_sc_hd__buf_1
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08363_ input27/X _08363_/B VGND VGND VPWR VPWR _08364_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08294_ _08311_/A input21/X _08312_/A _08314_/A VGND VGND VPWR VPWR _08309_/A sky130_fd_sc_hd__o22a_1
XFILLER_3_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09817_ _09817_/A _09817_/B _09826_/B VGND VGND VPWR VPWR _09818_/B sky130_fd_sc_hd__or3_1
XFILLER_46_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09748_ _09750_/B VGND VGND VPWR VPWR _10034_/A sky130_fd_sc_hd__inv_2
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11710_ _11710_/A VGND VGND VPWR VPWR _11771_/A sky130_fd_sc_hd__inv_2
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09679_ _08667_/A _09681_/B _09799_/B VGND VGND VPWR VPWR _09829_/B sky130_fd_sc_hd__o21ai_2
XFILLER_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12690_/A _12690_/B VGND VGND VPWR VPWR _12690_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _12452_/A _11641_/B VGND VGND VPWR VPWR _11641_/X sky130_fd_sc_hd__or2_1
X_14360_ _15948_/A VGND VGND VPWR VPWR _14378_/B sky130_fd_sc_hd__inv_2
X_11572_ _12404_/A VGND VGND VPWR VPWR _15437_/A sky130_fd_sc_hd__buf_1
X_13311_ _14858_/A _13306_/B _13306_/Y VGND VGND VPWR VPWR _13311_/Y sky130_fd_sc_hd__o21ai_1
X_10523_ _11833_/A _10523_/B VGND VGND VPWR VPWR _10523_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 wbs_dat_i[10] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__buf_1
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14291_ _15982_/A _14405_/B VGND VGND VPWR VPWR _14291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16030_ _16030_/A _16030_/B VGND VGND VPWR VPWR _16030_/Y sky130_fd_sc_hd__nand2_1
X_13242_ _14439_/A VGND VGND VPWR VPWR _14733_/A sky130_fd_sc_hd__buf_1
X_10454_ _10453_/Y _10370_/X _10379_/Y VGND VGND VPWR VPWR _10454_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13173_ _13104_/X _13172_/Y _13104_/X _13172_/Y VGND VGND VPWR VPWR _13186_/B sky130_fd_sc_hd__a2bb2o_1
X_10385_ _10251_/A _10384_/Y _10251_/Y _10384_/A _10472_/A VGND VGND VPWR VPWR _11803_/A
+ sky130_fd_sc_hd__o221a_2
X_12124_ _12052_/X _12123_/Y _12052_/X _12123_/Y VGND VGND VPWR VPWR _12141_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12055_ _12055_/A _12055_/B VGND VGND VPWR VPWR _12055_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11006_ _13898_/A _11093_/B VGND VGND VPWR VPWR _11186_/A sky130_fd_sc_hd__and2_1
XFILLER_38_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15814_ _15737_/Y _15812_/X _15813_/Y VGND VGND VPWR VPWR _15814_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15745_ _14915_/X _15744_/X _14915_/X _15744_/X VGND VGND VPWR VPWR _15746_/B sky130_fd_sc_hd__a2bb2oi_1
X_12957_ _14836_/A _13034_/B VGND VGND VPWR VPWR _13039_/A sky130_fd_sc_hd__and2_1
XFILLER_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15676_ _15622_/Y _15674_/X _15675_/Y VGND VGND VPWR VPWR _15676_/X sky130_fd_sc_hd__o21a_1
X_11908_ _11870_/Y _11906_/Y _11907_/Y VGND VGND VPWR VPWR _11979_/A sky130_fd_sc_hd__o21ai_1
X_12888_ _12934_/A VGND VGND VPWR VPWR _14469_/A sky130_fd_sc_hd__buf_1
XFILLER_61_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14627_ _14627_/A VGND VGND VPWR VPWR _15337_/A sky130_fd_sc_hd__buf_1
X_11839_ _11839_/A _11839_/B VGND VGND VPWR VPWR _11839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14558_ _14513_/X _14557_/X _14513_/X _14557_/X VGND VGND VPWR VPWR _14578_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14489_ _14489_/A VGND VGND VPWR VPWR _15202_/A sky130_fd_sc_hd__buf_1
X_13509_ _10830_/X _13488_/X _10830_/X _13488_/X VGND VGND VPWR VPWR _13510_/B sky130_fd_sc_hd__o2bb2a_1
X_16228_ _16228_/A VGND VGND VPWR VPWR _16228_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16159_ _15816_/X _16158_/X _15816_/X _16158_/X VGND VGND VPWR VPWR _16160_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08981_ _08885_/X _08979_/X _11357_/B VGND VGND VPWR VPWR _08981_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09602_ _09552_/X _09601_/Y _09552_/X _09601_/Y VGND VGND VPWR VPWR _09656_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09533_ _09555_/A _09555_/B VGND VGND VPWR VPWR _09595_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09464_ _10017_/A _08623_/A _09457_/Y _09463_/X VGND VGND VPWR VPWR _09464_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09395_ _11128_/A VGND VGND VPWR VPWR _09396_/A sky130_fd_sc_hd__buf_1
X_08415_ _08414_/A _08348_/Y _08414_/Y _08348_/A _08419_/A VGND VGND VPWR VPWR _09221_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08346_ input29/X _08346_/B VGND VGND VPWR VPWR _08347_/B sky130_fd_sc_hd__nor2_1
X_08277_ input25/X VGND VGND VPWR VPWR _08278_/A sky130_fd_sc_hd__inv_2
XFILLER_20_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10170_ _10251_/A _10170_/B VGND VGND VPWR VPWR _10170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13860_ _14745_/A _13860_/B VGND VGND VPWR VPWR _13860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13791_ _13864_/A _13790_/Y _13864_/A _13790_/Y VGND VGND VPWR VPWR _13793_/B sky130_fd_sc_hd__a2bb2o_1
X_12811_ _12771_/A _12771_/B _12771_/Y VGND VGND VPWR VPWR _12811_/Y sky130_fd_sc_hd__o21ai_1
X_15530_ _15526_/Y _15624_/A _15529_/Y VGND VGND VPWR VPWR _15534_/B sky130_fd_sc_hd__o21ai_2
XFILLER_103_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12694_/A _12694_/B _12694_/Y VGND VGND VPWR VPWR _12742_/X sky130_fd_sc_hd__a21o_1
X_15461_ _15461_/A _15461_/B VGND VGND VPWR VPWR _15461_/Y sky130_fd_sc_hd__nand2_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _11314_/Y _12672_/Y _11150_/Y VGND VGND VPWR VPWR _12674_/A sky130_fd_sc_hd__o21ai_1
X_14412_ _14412_/A VGND VGND VPWR VPWR _15193_/A sky130_fd_sc_hd__buf_1
XFILLER_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _12410_/A _11624_/B VGND VGND VPWR VPWR _11624_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15392_ _15392_/A _15398_/B VGND VGND VPWR VPWR _15468_/A sky130_fd_sc_hd__and2_1
X_14343_ _15875_/A _14257_/B _14257_/Y VGND VGND VPWR VPWR _14343_/Y sky130_fd_sc_hd__o21ai_1
X_11555_ _11555_/A _11554_/X VGND VGND VPWR VPWR _11555_/X sky130_fd_sc_hd__or2b_1
XFILLER_116_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14274_ _14274_/A VGND VGND VPWR VPWR _14274_/Y sky130_fd_sc_hd__inv_2
X_11486_ _13042_/A _11344_/B _11344_/Y _11283_/X VGND VGND VPWR VPWR _11486_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10506_ _13606_/A _10527_/B VGND VGND VPWR VPWR _10506_/Y sky130_fd_sc_hd__nor2_1
X_16013_ _16038_/A _16038_/B VGND VGND VPWR VPWR _16013_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13225_ _14741_/A _13300_/B VGND VGND VPWR VPWR _13225_/Y sky130_fd_sc_hd__nor2_1
X_10437_ _09313_/A _09313_/B _09313_/Y VGND VGND VPWR VPWR _10439_/A sky130_fd_sc_hd__o21ai_1
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13156_ _13198_/A _13198_/B VGND VGND VPWR VPWR _13156_/Y sky130_fd_sc_hd__nor2_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _10365_/Y _12700_/A _10299_/X _10367_/Y VGND VGND VPWR VPWR _10368_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12107_ _13898_/A _12153_/B VGND VGND VPWR VPWR _12204_/A sky130_fd_sc_hd__and2_1
X_13087_ _15261_/A _13107_/B VGND VGND VPWR VPWR _13087_/Y sky130_fd_sc_hd__nor2_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10296_/A _10325_/B _10295_/X _10298_/Y VGND VGND VPWR VPWR _10299_/X sky130_fd_sc_hd__o22a_1
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12038_ _12038_/A _11964_/X VGND VGND VPWR VPWR _12038_/X sky130_fd_sc_hd__or2b_1
XFILLER_78_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13989_ _13989_/A _13989_/B VGND VGND VPWR VPWR _13989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15728_ _15728_/A _15728_/B VGND VGND VPWR VPWR _16114_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15659_ _12610_/A _15658_/A _12610_/Y _15658_/Y _15655_/B VGND VGND VPWR VPWR _16027_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_61_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09180_ _09431_/A _09180_/B VGND VGND VPWR VPWR _09180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08964_ _08963_/Y _08859_/X _08963_/Y _08859_/X VGND VGND VPWR VPWR _08968_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08895_ _08894_/Y _08863_/X _08894_/Y _08863_/X VGND VGND VPWR VPWR _08976_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09516_ _09484_/A _09484_/B _09484_/Y _09515_/X VGND VGND VPWR VPWR _09516_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _12063_/A VGND VGND VPWR VPWR _10921_/A sky130_fd_sc_hd__inv_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09378_ _09472_/B _09860_/A _09353_/A VGND VGND VPWR VPWR _09378_/X sky130_fd_sc_hd__o21a_1
X_08329_ _08329_/A VGND VGND VPWR VPWR _08329_/Y sky130_fd_sc_hd__inv_2
X_11340_ _11296_/X _11339_/Y _11296_/X _11339_/Y VGND VGND VPWR VPWR _11491_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13010_ _13677_/A _13010_/B VGND VGND VPWR VPWR _13010_/Y sky130_fd_sc_hd__nand2_1
X_11271_ _11504_/A VGND VGND VPWR VPWR _13786_/A sky130_fd_sc_hd__buf_1
XFILLER_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10222_ _10222_/A VGND VGND VPWR VPWR _10222_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10153_ _10155_/A VGND VGND VPWR VPWR _10242_/B sky130_fd_sc_hd__buf_1
XFILLER_121_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14961_ _14971_/A _14971_/B VGND VGND VPWR VPWR _14961_/Y sky130_fd_sc_hd__nand2_1
X_10084_ _10043_/X _10082_/X _11142_/B VGND VGND VPWR VPWR _10084_/X sky130_fd_sc_hd__o21a_1
X_14892_ _15529_/A _14912_/B VGND VGND VPWR VPWR _14892_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13912_ _13849_/X _13911_/Y _13849_/X _13911_/Y VGND VGND VPWR VPWR _13950_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13843_ _13828_/Y _13841_/X _13842_/Y VGND VGND VPWR VPWR _13843_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15513_ _15470_/A _15470_/B _15470_/Y VGND VGND VPWR VPWR _15513_/Y sky130_fd_sc_hd__o21ai_1
X_13774_ _13804_/A _13772_/X _13773_/X VGND VGND VPWR VPWR _13774_/X sky130_fd_sc_hd__o21a_1
X_10986_ _11138_/A _12688_/A _10985_/Y VGND VGND VPWR VPWR _10986_/X sky130_fd_sc_hd__a21o_1
X_12725_ _12719_/X _12724_/X _12719_/X _12724_/X VGND VGND VPWR VPWR _12785_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15444_ _15444_/A _15414_/X VGND VGND VPWR VPWR _15444_/X sky130_fd_sc_hd__or2b_1
X_12656_ _10282_/Y _10206_/A _10349_/A VGND VGND VPWR VPWR _12656_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12587_ _12587_/A VGND VGND VPWR VPWR _12587_/Y sky130_fd_sc_hd__inv_2
X_15375_ _15375_/A _15341_/X VGND VGND VPWR VPWR _15375_/X sky130_fd_sc_hd__or2b_1
X_11607_ _11607_/A VGND VGND VPWR VPWR _11607_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14326_ _14265_/A _14325_/Y _14326_/B1 _14325_/Y VGND VGND VPWR VPWR _14388_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11538_ _13496_/A _11626_/B _13496_/A _11626_/B VGND VGND VPWR VPWR _11538_/X sky130_fd_sc_hd__a2bb2o_1
X_14257_ _15875_/A _14257_/B VGND VGND VPWR VPWR _14257_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11469_ _09184_/Y _11468_/A _09184_/A _11468_/Y _09204_/X VGND VGND VPWR VPWR _13313_/A
+ sky130_fd_sc_hd__a221o_4
X_14188_ _14116_/X _14187_/Y _14116_/X _14187_/Y VGND VGND VPWR VPWR _14189_/B sky130_fd_sc_hd__a2bb2oi_1
X_13208_ _13140_/X _13207_/X _13140_/X _13207_/X VGND VGND VPWR VPWR _13452_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13139_ _13139_/A _13139_/B VGND VGND VPWR VPWR _13139_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08680_ _08679_/A _08679_/B _08678_/Y _08679_/X VGND VGND VPWR VPWR _08680_/X sky130_fd_sc_hd__o22a_2
XFILLER_66_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09301_ _09301_/A VGND VGND VPWR VPWR _09301_/Y sky130_fd_sc_hd__inv_2
X_09232_ _09232_/A _09232_/B VGND VGND VPWR VPWR _09678_/A sky130_fd_sc_hd__or2_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09163_ _08757_/Y _09160_/A _08757_/A _09160_/Y VGND VGND VPWR VPWR _10009_/B sky130_fd_sc_hd__o22a_1
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09094_ _09705_/A VGND VGND VPWR VPWR _09415_/A sky130_fd_sc_hd__buf_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09996_ _09965_/X _11307_/A _11306_/B VGND VGND VPWR VPWR _11510_/A sky130_fd_sc_hd__o21a_1
X_08947_ _08946_/Y _08857_/X _08946_/Y _08857_/X VGND VGND VPWR VPWR _08952_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_57_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08878_ _08770_/A _08770_/B _08770_/Y VGND VGND VPWR VPWR _08878_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10840_ _13701_/A _10935_/B _10839_/Y VGND VGND VPWR VPWR _10840_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10771_ _13088_/A _10747_/B _10747_/Y _10770_/X VGND VGND VPWR VPWR _10771_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12510_ _12509_/A _12509_/B _12509_/Y _12501_/X VGND VGND VPWR VPWR _12637_/B sky130_fd_sc_hd__o211a_1
XFILLER_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13490_ _11136_/Y _12087_/A _10985_/Y _13489_/X VGND VGND VPWR VPWR _13490_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12441_ _13872_/A _12440_/B _12440_/X _12368_/X VGND VGND VPWR VPWR _12441_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12372_ _13496_/A VGND VGND VPWR VPWR _12435_/A sky130_fd_sc_hd__inv_2
X_15160_ _12380_/A _15101_/X _12379_/X VGND VGND VPWR VPWR _15161_/A sky130_fd_sc_hd__o21ai_1
XFILLER_125_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14111_ _14054_/X _14110_/X _14054_/X _14110_/X VGND VGND VPWR VPWR _14111_/Y sky130_fd_sc_hd__a2bb2oi_1
X_15091_ _15078_/A _15078_/B _15078_/Y _15090_/X VGND VGND VPWR VPWR _15091_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11323_ _11322_/A _11321_/Y _11322_/Y _11321_/A _11526_/A VGND VGND VPWR VPWR _11518_/B
+ sky130_fd_sc_hd__a221o_1
X_11254_ _14036_/A _11230_/B _11230_/Y _11253_/X VGND VGND VPWR VPWR _11254_/X sky130_fd_sc_hd__a2bb2o_1
X_14042_ _13939_/X _14041_/X _13939_/X _14041_/X VGND VGND VPWR VPWR _14043_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10205_ _10346_/B _10899_/B VGND VGND VPWR VPWR _10206_/A sky130_fd_sc_hd__or2_1
X_11185_ _14060_/A VGND VGND VPWR VPWR _15446_/A sky130_fd_sc_hd__buf_1
X_15993_ _15993_/A _15972_/X VGND VGND VPWR VPWR _15993_/X sky130_fd_sc_hd__or2b_1
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10136_ _10120_/A _10120_/B _10120_/X VGND VGND VPWR VPWR _10139_/A sky130_fd_sc_hd__a21bo_1
XFILLER_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14944_ _14944_/A _14944_/B VGND VGND VPWR VPWR _14944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10067_ _10067_/A _10067_/B VGND VGND VPWR VPWR _10067_/X sky130_fd_sc_hd__or2_1
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14875_ _15546_/A _14922_/B VGND VGND VPWR VPWR _14875_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13826_ _13826_/A _13759_/X VGND VGND VPWR VPWR _13826_/X sky130_fd_sc_hd__or2b_1
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13757_ _13757_/A _13757_/B VGND VGND VPWR VPWR _13757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10969_ _11604_/A _10969_/B VGND VGND VPWR VPWR _10970_/A sky130_fd_sc_hd__or2_1
X_12708_ _13479_/A _12707_/X _10289_/X VGND VGND VPWR VPWR _12708_/X sky130_fd_sc_hd__o21a_1
X_13688_ _13680_/Y _13686_/Y _13687_/Y VGND VGND VPWR VPWR _13688_/X sky130_fd_sc_hd__o21a_1
X_15427_ _12428_/A _15163_/B _15163_/Y _15165_/Y VGND VGND VPWR VPWR _15427_/Y sky130_fd_sc_hd__o2bb2ai_1
X_12639_ _12639_/A _12639_/B VGND VGND VPWR VPWR _12639_/X sky130_fd_sc_hd__or2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15358_ _15352_/X _15357_/X _15352_/X _15357_/X VGND VGND VPWR VPWR _15420_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14309_ _14309_/A _14309_/B VGND VGND VPWR VPWR _15964_/A sky130_fd_sc_hd__or2_1
X_15289_ _15289_/A _15289_/B VGND VGND VPWR VPWR _15289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09850_ _09848_/A _09848_/B _09849_/Y VGND VGND VPWR VPWR _09850_/Y sky130_fd_sc_hd__o21ai_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08801_ _08801_/A VGND VGND VPWR VPWR _10128_/A sky130_fd_sc_hd__inv_2
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09782_/A _09782_/B VGND VGND VPWR VPWR _09781_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08732_ _08713_/A _08713_/B _08713_/X _08731_/Y VGND VGND VPWR VPWR _08733_/A sky130_fd_sc_hd__a22o_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08663_ _09677_/A _08663_/B VGND VGND VPWR VPWR _08665_/A sky130_fd_sc_hd__or2_1
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _09455_/B VGND VGND VPWR VPWR _08715_/B sky130_fd_sc_hd__inv_2
XFILLER_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09215_ _09551_/A _09728_/A VGND VGND VPWR VPWR _09216_/A sky130_fd_sc_hd__or2_1
XFILLER_108_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09146_ _09146_/A VGND VGND VPWR VPWR _09146_/X sky130_fd_sc_hd__buf_1
XFILLER_108_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09077_ _10012_/B _09077_/B VGND VGND VPWR VPWR _09078_/B sky130_fd_sc_hd__or2_1
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09979_ _09970_/Y _09977_/Y _09978_/Y VGND VGND VPWR VPWR _09981_/B sky130_fd_sc_hd__o21ai_1
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12990_ _12990_/A VGND VGND VPWR VPWR _13015_/A sky130_fd_sc_hd__inv_2
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11941_ _11906_/A _11940_/Y _11906_/A _11940_/Y VGND VGND VPWR VPWR _11974_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14660_ _15345_/A _14660_/B VGND VGND VPWR VPWR _14660_/Y sky130_fd_sc_hd__nand2_1
X_11872_ _11842_/X _11871_/Y _11842_/X _11871_/Y VGND VGND VPWR VPWR _11904_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14591_ _14523_/X _14537_/A _14536_/X VGND VGND VPWR VPWR _14591_/X sky130_fd_sc_hd__o21a_1
X_13611_ _12916_/Y _12917_/X _12916_/A _12915_/Y VGND VGND VPWR VPWR _13612_/A sky130_fd_sc_hd__a22o_1
XFILLER_60_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10823_ _10823_/A VGND VGND VPWR VPWR _10823_/Y sky130_fd_sc_hd__inv_2
X_16330_ _16330_/A _16330_/B VGND VGND VPWR VPWR _16330_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13542_ _15051_/A _13501_/B _13501_/Y _13541_/X VGND VGND VPWR VPWR _13542_/X sky130_fd_sc_hd__a2bb2o_1
X_10754_ _10627_/X _10753_/Y _10627_/X _10753_/Y VGND VGND VPWR VPWR _10769_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16261_ _16194_/Y _16259_/X _16260_/Y VGND VGND VPWR VPWR _16261_/X sky130_fd_sc_hd__o21a_1
X_13473_ _14368_/A VGND VGND VPWR VPWR _14353_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10685_ _10685_/A VGND VGND VPWR VPWR _10685_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16192_ _16192_/A _16192_/B VGND VGND VPWR VPWR _16260_/B sky130_fd_sc_hd__or2_1
X_15212_ _15212_/A _15212_/B VGND VGND VPWR VPWR _15212_/X sky130_fd_sc_hd__or2_1
X_12424_ _11609_/A _11691_/B _12422_/Y _12423_/Y VGND VGND VPWR VPWR _12424_/X sky130_fd_sc_hd__o22a_2
X_12355_ _12300_/A _12300_/B _12300_/Y _12509_/A VGND VGND VPWR VPWR _12409_/A sky130_fd_sc_hd__a2bb2o_1
X_15143_ _15143_/A _15143_/B VGND VGND VPWR VPWR _15143_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11306_ _09965_/X _11306_/B VGND VGND VPWR VPWR _11307_/B sky130_fd_sc_hd__and2b_1
X_12286_ _12363_/A _12285_/Y _12363_/A _12285_/Y VGND VGND VPWR VPWR _12360_/B sky130_fd_sc_hd__a2bb2o_1
X_15074_ _15033_/X _15073_/X _15033_/X _15073_/X VGND VGND VPWR VPWR _15075_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14025_ _14028_/A VGND VGND VPWR VPWR _15458_/A sky130_fd_sc_hd__buf_1
X_11237_ _11237_/A _11249_/B VGND VGND VPWR VPWR _14043_/A sky130_fd_sc_hd__or2_1
XFILLER_122_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11168_ _13720_/A _11288_/B _11167_/Y VGND VGND VPWR VPWR _11168_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10119_ _10119_/A _10119_/B VGND VGND VPWR VPWR _10120_/A sky130_fd_sc_hd__or2_1
X_15976_ _15984_/A _15984_/B VGND VGND VPWR VPWR _15976_/Y sky130_fd_sc_hd__nand2_1
X_11099_ _12259_/A VGND VGND VPWR VPWR _13713_/A sky130_fd_sc_hd__buf_1
XFILLER_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14927_ _14867_/Y _14925_/X _14926_/Y VGND VGND VPWR VPWR _14927_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14858_ _14858_/A _14858_/B VGND VGND VPWR VPWR _14858_/X sky130_fd_sc_hd__or2_1
XFILLER_90_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13809_ _14611_/A _13854_/B VGND VGND VPWR VPWR _13809_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14789_ _14734_/X _14788_/X _14734_/X _14788_/X VGND VGND VPWR VPWR _14790_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16459_ _08229_/A _16459_/D VGND VGND VPWR VPWR _16459_/Q sky130_fd_sc_hd__dfxtp_1
X_09000_ _11391_/A VGND VGND VPWR VPWR _11569_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09902_ _09903_/A _09903_/B VGND VGND VPWR VPWR _10654_/B sky130_fd_sc_hd__and2_1
X_09833_ _09833_/A VGND VGND VPWR VPWR _09833_/Y sky130_fd_sc_hd__inv_2
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09733_/A _09733_/B _09736_/A VGND VGND VPWR VPWR _10049_/A sky130_fd_sc_hd__a21bo_1
XFILLER_82_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08715_ _08715_/A _08715_/B VGND VGND VPWR VPWR _08715_/X sky130_fd_sc_hd__or2_1
X_09695_ _09695_/A _09695_/B VGND VGND VPWR VPWR _09698_/A sky130_fd_sc_hd__or2_1
Xrebuffer20 rebuffer21/X VGND VGND VPWR VPWR rebuffer20/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer31 _16313_/A2 VGND VGND VPWR VPWR _16316_/A sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08646_ _08645_/X _08407_/Y _08645_/X _08407_/Y VGND VGND VPWR VPWR _08647_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_27_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _09454_/B VGND VGND VPWR VPWR _09553_/A sky130_fd_sc_hd__buf_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10470_ _09313_/A _10254_/B _10255_/A VGND VGND VPWR VPWR _10471_/A sky130_fd_sc_hd__o21ai_1
X_09129_ _09553_/B _09035_/B _09036_/B VGND VGND VPWR VPWR _09130_/A sky130_fd_sc_hd__a21bo_1
X_12140_ _12225_/A _12138_/X _12139_/X VGND VGND VPWR VPWR _12140_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12071_ _13641_/A _12071_/B VGND VGND VPWR VPWR _12071_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11022_ _13552_/A VGND VGND VPWR VPWR _12848_/A sky130_fd_sc_hd__buf_1
X_15830_ _14407_/Y _15829_/X _14407_/Y _15829_/X VGND VGND VPWR VPWR _16238_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_49_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15761_ _14909_/X _15760_/X _14909_/X _15760_/X VGND VGND VPWR VPWR _15762_/B sky130_fd_sc_hd__a2bb2oi_1
X_12973_ _14524_/A _13026_/B VGND VGND VPWR VPWR _13060_/A sky130_fd_sc_hd__and2_1
XFILLER_64_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15692_ _15700_/A _15692_/B VGND VGND VPWR VPWR _16053_/A sky130_fd_sc_hd__or2_1
X_14712_ _15333_/A _14648_/B _14648_/Y VGND VGND VPWR VPWR _14712_/Y sky130_fd_sc_hd__o21ai_1
X_11924_ _11925_/A _11925_/B VGND VGND VPWR VPWR _11926_/A sky130_fd_sc_hd__and2_1
X_14643_ _13096_/X _14642_/Y _13096_/X _14642_/Y VGND VGND VPWR VPWR _14644_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11855_ _10459_/A _11807_/A _10554_/B _11854_/Y VGND VGND VPWR VPWR _11856_/A sky130_fd_sc_hd__o22a_1
X_14574_ _15272_/A _14574_/B VGND VGND VPWR VPWR _14574_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11786_ _11719_/B _11785_/X _11719_/B _11785_/X VGND VGND VPWR VPWR _11787_/B sky130_fd_sc_hd__a2bb2o_1
X_10806_ _11988_/A VGND VGND VPWR VPWR _13510_/A sky130_fd_sc_hd__buf_1
XFILLER_13_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16313_ _16249_/A _16313_/A2 _16249_/Y VGND VGND VPWR VPWR _16313_/Y sky130_fd_sc_hd__o21ai_1
X_10737_ _10634_/A _10736_/Y _10634_/A _10736_/Y VGND VGND VPWR VPWR _10738_/B sky130_fd_sc_hd__a2bb2o_1
X_13525_ _13525_/A _13525_/B VGND VGND VPWR VPWR _13525_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16244_ _16244_/A VGND VGND VPWR VPWR _16457_/S sky130_fd_sc_hd__buf_1
XFILLER_127_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13456_ _13454_/X _13455_/Y _13454_/X _13455_/Y VGND VGND VPWR VPWR _13456_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12407_ _12407_/A _12407_/B VGND VGND VPWR VPWR _12407_/Y sky130_fd_sc_hd__nand2_1
X_10668_ _11916_/A VGND VGND VPWR VPWR _13513_/A sky130_fd_sc_hd__buf_1
XFILLER_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16175_ _15812_/X _16174_/X _15812_/X _16174_/X VGND VGND VPWR VPWR _16176_/B sky130_fd_sc_hd__a2bb2o_1
X_13387_ _14126_/A _13442_/B VGND VGND VPWR VPWR _13387_/Y sky130_fd_sc_hd__nor2_1
X_10599_ _10528_/X _10598_/Y _10528_/X _10598_/Y VGND VGND VPWR VPWR _10635_/B sky130_fd_sc_hd__a2bb2o_1
X_12338_ _12240_/X _12337_/Y _12240_/X _12337_/Y VGND VGND VPWR VPWR _12569_/A sky130_fd_sc_hd__a2bb2o_1
X_15126_ _15069_/A _15069_/B _15069_/Y VGND VGND VPWR VPWR _15126_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15057_ _15057_/A _15057_/B VGND VGND VPWR VPWR _15057_/Y sky130_fd_sc_hd__nand2_1
X_12269_ _11145_/A _12176_/A _11314_/B _12268_/Y VGND VGND VPWR VPWR _12270_/A sky130_fd_sc_hd__o22a_1
X_14008_ _13959_/X _14007_/Y _13959_/X _14007_/Y VGND VGND VPWR VPWR _14064_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15959_ _16008_/A _15957_/X _15958_/X VGND VGND VPWR VPWR _15959_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08500_ _08589_/A VGND VGND VPWR VPWR _08701_/A sky130_fd_sc_hd__buf_1
X_09480_ _08749_/A _09520_/S _08749_/A _09520_/S VGND VGND VPWR VPWR _09518_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08431_ _09209_/A VGND VGND VPWR VPWR _08713_/A sky130_fd_sc_hd__inv_2
XFILLER_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08362_ _08275_/A input10/X _08387_/B _08361_/Y VGND VGND VPWR VPWR _08366_/A sky130_fd_sc_hd__o22a_1
X_08293_ _08316_/A input20/X _08317_/A _08319_/A VGND VGND VPWR VPWR _08314_/A sky130_fd_sc_hd__o22a_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09816_ _09809_/X _08839_/Y _09809_/X _08839_/Y VGND VGND VPWR VPWR _09818_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09747_ _09791_/A _09791_/B _09791_/A _09791_/B VGND VGND VPWR VPWR _09750_/B sky130_fd_sc_hd__a2bb2o_2
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09678_ _09678_/A _09680_/A VGND VGND VPWR VPWR _09799_/B sky130_fd_sc_hd__or2_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08629_ _09458_/B VGND VGND VPWR VPWR _09538_/A sky130_fd_sc_hd__buf_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11640_ _11637_/X _11639_/X _11637_/X _11639_/X VGND VGND VPWR VPWR _11641_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11571_ _12494_/A VGND VGND VPWR VPWR _15554_/A sky130_fd_sc_hd__buf_1
X_13310_ _14068_/A _13309_/B _13309_/Y VGND VGND VPWR VPWR _13310_/X sky130_fd_sc_hd__a21o_1
X_10522_ _10522_/A VGND VGND VPWR VPWR _10522_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14290_ _14167_/X _14289_/X _14167_/X _14289_/X VGND VGND VPWR VPWR _14405_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13241_ _15069_/A VGND VGND VPWR VPWR _14439_/A sky130_fd_sc_hd__inv_2
X_10453_ _11805_/A _10453_/B VGND VGND VPWR VPWR _10453_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13172_ _15264_/A _13105_/B _13105_/Y VGND VGND VPWR VPWR _13172_/Y sky130_fd_sc_hd__o21ai_1
X_10384_ _10384_/A VGND VGND VPWR VPWR _10384_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12123_ _13188_/A _12053_/B _12053_/Y VGND VGND VPWR VPWR _12123_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12054_ _12034_/Y _12052_/X _12053_/Y VGND VGND VPWR VPWR _12054_/X sky130_fd_sc_hd__o21a_1
X_11005_ _10923_/X _11004_/X _10923_/X _11004_/X VGND VGND VPWR VPWR _11093_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15813_ _16112_/A _15813_/B VGND VGND VPWR VPWR _15813_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15744_ _14916_/A _14916_/B _14916_/Y VGND VGND VPWR VPWR _15744_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12956_ _12945_/X _12955_/Y _12945_/X _12955_/Y VGND VGND VPWR VPWR _13034_/B sky130_fd_sc_hd__a2bb2o_1
X_15675_ _15675_/A _15675_/B VGND VGND VPWR VPWR _15675_/Y sky130_fd_sc_hd__nand2_1
X_11907_ _11907_/A _11907_/B VGND VGND VPWR VPWR _11907_/Y sky130_fd_sc_hd__nand2_1
X_12887_ _14477_/A _12936_/B VGND VGND VPWR VPWR _12887_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _15339_/A _14654_/B VGND VGND VPWR VPWR _14626_/Y sky130_fd_sc_hd__nor2_1
X_11838_ _11827_/Y _11836_/X _11837_/Y VGND VGND VPWR VPWR _11838_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/A _14514_/X VGND VGND VPWR VPWR _14557_/X sky130_fd_sc_hd__or2b_1
XFILLER_119_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11769_ _11798_/B _11768_/Y _11798_/B _11768_/Y VGND VGND VPWR VPWR _11770_/B sky130_fd_sc_hd__o2bb2a_1
X_13508_ _13510_/A VGND VGND VPWR VPWR _15042_/A sky130_fd_sc_hd__buf_1
X_14488_ _15199_/A _14518_/B VGND VGND VPWR VPWR _14549_/A sky130_fd_sc_hd__and2_1
X_16227_ _16227_/A VGND VGND VPWR VPWR _16227_/Y sky130_fd_sc_hd__inv_2
X_13439_ _13393_/Y _13437_/X _13438_/Y VGND VGND VPWR VPWR _13439_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16158_ _15817_/A _15817_/B _15817_/Y VGND VGND VPWR VPWR _16158_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15109_ _15099_/X _15108_/Y _15099_/X _15108_/Y VGND VGND VPWR VPWR _15110_/B sky130_fd_sc_hd__a2bb2o_1
X_16089_ _16089_/A _16089_/B VGND VGND VPWR VPWR _16089_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08980_ _08980_/A _08980_/B VGND VGND VPWR VPWR _11357_/B sky130_fd_sc_hd__or2_1
XFILLER_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09601_ _09601_/A _09601_/B VGND VGND VPWR VPWR _09601_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09532_ _09532_/A VGND VGND VPWR VPWR _09532_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09463_ _09458_/Y _09461_/X _09462_/X VGND VGND VPWR VPWR _09463_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08414_ _08414_/A VGND VGND VPWR VPWR _08414_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09394_ _09330_/A _09330_/B _09330_/Y _09393_/X VGND VGND VPWR VPWR _11128_/A sky130_fd_sc_hd__o211a_1
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08345_ _08343_/Y _08344_/A _08343_/A _08344_/Y _08304_/A VGND VGND VPWR VPWR _09217_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08276_ input9/X VGND VGND VPWR VPWR _08276_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12810_ _12848_/A _12848_/B VGND VGND VPWR VPWR _12810_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13790_ _15113_/A _13865_/B _13789_/Y VGND VGND VPWR VPWR _13790_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12741_ _12775_/A _12775_/B VGND VGND VPWR VPWR _12741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15460_ _15403_/X _15459_/X _15403_/X _15459_/X VGND VGND VPWR VPWR _15461_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12672_ _12672_/A VGND VGND VPWR VPWR _12672_/Y sky130_fd_sc_hd__inv_2
X_14411_ _15246_/A VGND VGND VPWR VPWR _14588_/A sky130_fd_sc_hd__buf_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A VGND VGND VPWR VPWR _11624_/B sky130_fd_sc_hd__inv_2
X_15391_ _15330_/X _15390_/Y _15330_/X _15390_/Y VGND VGND VPWR VPWR _15398_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14342_ _14384_/A _15954_/A VGND VGND VPWR VPWR _15628_/A sky130_fd_sc_hd__and2_1
X_11554_ _14832_/A _11554_/B VGND VGND VPWR VPWR _11554_/X sky130_fd_sc_hd__or2_1
XFILLER_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14273_ _14192_/Y _14271_/Y _14272_/Y VGND VGND VPWR VPWR _14274_/A sky130_fd_sc_hd__o21ai_2
X_11485_ _13206_/A VGND VGND VPWR VPWR _12397_/A sky130_fd_sc_hd__inv_2
X_10505_ _10433_/X _10504_/X _10433_/X _10504_/X VGND VGND VPWR VPWR _10527_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16012_ _15955_/X _16011_/X _15955_/X _16011_/X VGND VGND VPWR VPWR _16038_/B sky130_fd_sc_hd__a2bb2o_1
X_13224_ _13201_/X _13223_/Y _13201_/X _13223_/Y VGND VGND VPWR VPWR _13300_/B sky130_fd_sc_hd__a2bb2o_1
X_10436_ _13560_/A _10392_/B _10392_/X _10435_/X VGND VGND VPWR VPWR _10436_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13155_ _13116_/X _13154_/Y _13116_/X _13154_/Y VGND VGND VPWR VPWR _13198_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10367_ _10367_/A _11750_/A VGND VGND VPWR VPWR _10367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12106_ _12064_/X _12105_/Y _12064_/X _12105_/Y VGND VGND VPWR VPWR _12153_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13086_ _13014_/X _13085_/X _13014_/X _13085_/X VGND VGND VPWR VPWR _13107_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10325_/A _12701_/A VGND VGND VPWR VPWR _10298_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12037_ _12037_/A _12051_/B VGND VGND VPWR VPWR _12037_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13988_ _13986_/X _13987_/X _13986_/X _13987_/X VGND VGND VPWR VPWR _13989_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15727_ _14921_/X _15726_/X _14921_/X _15726_/X VGND VGND VPWR VPWR _15728_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12939_ _12883_/Y _12937_/X _12938_/Y VGND VGND VPWR VPWR _12939_/X sky130_fd_sc_hd__o21a_1
X_15658_ _15658_/A VGND VGND VPWR VPWR _15658_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14609_ _14589_/X _14608_/Y _14589_/X _14608_/Y VGND VGND VPWR VPWR _14662_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15589_ _16046_/A VGND VGND VPWR VPWR _15683_/A sky130_fd_sc_hd__inv_2
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08963_ _08962_/X _10125_/A _08827_/Y VGND VGND VPWR VPWR _08963_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08894_ _08893_/X _08793_/B _08793_/Y VGND VGND VPWR VPWR _08894_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09515_ _09486_/A _09486_/B _09486_/Y _09514_/X VGND VGND VPWR VPWR _09515_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ _09248_/A _09428_/A _09263_/A _09428_/Y _10926_/A VGND VGND VPWR VPWR _12063_/A
+ sky130_fd_sc_hd__a221o_2
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09377_ _09431_/B _09377_/B VGND VGND VPWR VPWR _09377_/X sky130_fd_sc_hd__or2_1
X_08328_ _08328_/A VGND VGND VPWR VPWR _08328_/Y sky130_fd_sc_hd__inv_2
X_08259_ input31/X VGND VGND VPWR VPWR _08260_/B sky130_fd_sc_hd__inv_2
XFILLER_20_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11270_ _11269_/A _11269_/B _11269_/Y _09393_/X VGND VGND VPWR VPWR _11504_/A sky130_fd_sc_hd__o211a_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10221_ _10180_/A _10180_/B _10180_/Y VGND VGND VPWR VPWR _10222_/A sky130_fd_sc_hd__o21ai_1
XFILLER_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10152_ _10116_/A _10116_/B _10117_/A VGND VGND VPWR VPWR _10155_/A sky130_fd_sc_hd__a21bo_1
X_14960_ _14957_/X _14959_/X _14957_/X _14959_/X VGND VGND VPWR VPWR _14971_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10083_ _10083_/A _10083_/B VGND VGND VPWR VPWR _11142_/B sky130_fd_sc_hd__or2_1
X_13911_ _14619_/A _13850_/B _13850_/Y VGND VGND VPWR VPWR _13911_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14891_ _14819_/X _14890_/X _14819_/X _14890_/X VGND VGND VPWR VPWR _14912_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13842_ _14635_/A _13842_/B VGND VGND VPWR VPWR _13842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13773_ _13773_/A _13773_/B VGND VGND VPWR VPWR _13773_/X sky130_fd_sc_hd__or2_1
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15512_ _15512_/A _15512_/B VGND VGND VPWR VPWR _15512_/X sky130_fd_sc_hd__and2_1
X_12724_ _12682_/A _12682_/B _12682_/Y VGND VGND VPWR VPWR _12724_/X sky130_fd_sc_hd__a21o_1
X_10985_ _11138_/A _12172_/A VGND VGND VPWR VPWR _10985_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15443_ _15443_/A _15443_/B VGND VGND VPWR VPWR _15443_/X sky130_fd_sc_hd__and2_1
X_12655_ _12863_/A VGND VGND VPWR VPWR _15171_/A sky130_fd_sc_hd__buf_1
X_12586_ _12586_/A _11429_/X VGND VGND VPWR VPWR _12587_/A sky130_fd_sc_hd__or2b_1
X_15374_ _15410_/A _15410_/B VGND VGND VPWR VPWR _15450_/A sky130_fd_sc_hd__and2_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11606_ _10194_/A _11606_/A2 _10194_/Y VGND VGND VPWR VPWR _11607_/A sky130_fd_sc_hd__o21ai_1
X_14325_ _15866_/A _14266_/B _14266_/Y VGND VGND VPWR VPWR _14325_/Y sky130_fd_sc_hd__o21ai_1
X_11537_ _11517_/X _11536_/X _11517_/X _11536_/X VGND VGND VPWR VPWR _11626_/B sky130_fd_sc_hd__a2bb2o_1
X_14256_ _14256_/A VGND VGND VPWR VPWR _14256_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11468_ _11468_/A VGND VGND VPWR VPWR _11468_/Y sky130_fd_sc_hd__inv_2
X_14187_ _13440_/A _14121_/A _14119_/Y VGND VGND VPWR VPWR _14187_/Y sky130_fd_sc_hd__a21oi_1
X_13207_ _13144_/Y _13205_/X _13206_/Y VGND VGND VPWR VPWR _13207_/X sky130_fd_sc_hd__o21a_1
X_10419_ _10354_/X _10418_/Y _10354_/X _10418_/Y VGND VGND VPWR VPWR _10430_/B sky130_fd_sc_hd__a2bb2o_1
X_11399_ _11399_/A VGND VGND VPWR VPWR _11399_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13138_ _13126_/X _13137_/Y _13126_/X _13137_/Y VGND VGND VPWR VPWR _13139_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13069_ _13767_/A VGND VGND VPWR VPWR _15252_/A sky130_fd_sc_hd__buf_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09300_ _09298_/A _09298_/B _09297_/Y _09299_/Y VGND VGND VPWR VPWR _09304_/A sky130_fd_sc_hd__o22a_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09231_ _09540_/A _09684_/A VGND VGND VPWR VPWR _09231_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09162_ _08749_/Y _09161_/Y _08749_/Y _09161_/Y VGND VGND VPWR VPWR _10008_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09093_ _10017_/B _09072_/B _09073_/B VGND VGND VPWR VPWR _09705_/A sky130_fd_sc_hd__a21bo_1
XFILLER_89_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09995_ _09995_/A _09995_/B VGND VGND VPWR VPWR _11306_/B sky130_fd_sc_hd__or2_1
XFILLER_130_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08946_ _08946_/A VGND VGND VPWR VPWR _08946_/Y sky130_fd_sc_hd__inv_2
X_08877_ _08691_/X _08876_/Y _08691_/X _08876_/Y VGND VGND VPWR VPWR _08982_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10770_ _10896_/A _10767_/X _10769_/X VGND VGND VPWR VPWR _10770_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09429_ _09429_/A _09429_/B VGND VGND VPWR VPWR _09429_/X sky130_fd_sc_hd__or2_1
XFILLER_100_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12440_ _12440_/A _12440_/B VGND VGND VPWR VPWR _12440_/X sky130_fd_sc_hd__and2_1
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14110_ _15455_/A _14024_/B _14109_/A _14024_/B VGND VGND VPWR VPWR _14110_/X sky130_fd_sc_hd__a2bb2o_1
X_12371_ _12783_/A _12369_/B _12369_/X _12370_/Y VGND VGND VPWR VPWR _12435_/B sky130_fd_sc_hd__a22o_1
X_15090_ _15081_/A _15081_/B _15081_/Y _15089_/X VGND VGND VPWR VPWR _15090_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11322_ _11322_/A VGND VGND VPWR VPWR _11322_/Y sky130_fd_sc_hd__inv_2
X_11253_ _13341_/A _11236_/B _11236_/Y _11252_/X VGND VGND VPWR VPWR _11253_/X sky130_fd_sc_hd__a2bb2o_1
X_14041_ _14041_/A _13940_/X VGND VGND VPWR VPWR _14041_/X sky130_fd_sc_hd__or2b_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10204_ _08664_/X _09404_/Y _08671_/A _09403_/X VGND VGND VPWR VPWR _10899_/B sky130_fd_sc_hd__o22a_2
XFILLER_121_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11184_ _14015_/A VGND VGND VPWR VPWR _14060_/A sky130_fd_sc_hd__buf_1
XFILLER_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15992_ _15992_/A _15991_/X VGND VGND VPWR VPWR _15992_/X sky130_fd_sc_hd__or2b_1
XFILLER_67_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10135_ _10134_/A _10134_/B _10134_/X VGND VGND VPWR VPWR _10194_/A sky130_fd_sc_hd__a21bo_1
X_14943_ _15425_/A _14980_/B _14942_/Y VGND VGND VPWR VPWR _14943_/Y sky130_fd_sc_hd__o21ai_1
X_10066_ _10021_/X _10065_/Y _10021_/X _10065_/Y VGND VGND VPWR VPWR _10067_/B sky130_fd_sc_hd__a2bb2o_1
X_14874_ _14824_/X _14873_/X _14824_/X _14873_/X VGND VGND VPWR VPWR _14922_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13825_ _13825_/A VGND VGND VPWR VPWR _14635_/A sky130_fd_sc_hd__inv_2
XFILLER_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13756_ _13753_/A _13753_/B _13753_/Y _13755_/Y VGND VGND VPWR VPWR _13756_/X sky130_fd_sc_hd__o2bb2a_1
X_10968_ _10080_/X _10967_/X _10080_/X _10967_/X VGND VGND VPWR VPWR _10969_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13687_ _14501_/A _13687_/B VGND VGND VPWR VPWR _13687_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12707_ _10284_/Y _10350_/B _10206_/A _10349_/A VGND VGND VPWR VPWR _12707_/X sky130_fd_sc_hd__o22a_1
X_12638_ _14284_/A _12636_/X _12637_/X VGND VGND VPWR VPWR _12638_/X sky130_fd_sc_hd__o21a_1
X_10899_ _10904_/A _10899_/B VGND VGND VPWR VPWR _12047_/A sky130_fd_sc_hd__nand2b_1
X_15426_ _15159_/Y _15425_/Y _15171_/Y VGND VGND VPWR VPWR _15426_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ _12569_/A VGND VGND VPWR VPWR _12569_/Y sky130_fd_sc_hd__inv_2
X_15357_ _15357_/A _15353_/X VGND VGND VPWR VPWR _15357_/X sky130_fd_sc_hd__or2b_1
X_14308_ _13441_/X _14307_/X _13441_/X _14307_/X VGND VGND VPWR VPWR _14309_/B sky130_fd_sc_hd__a2bb2oi_1
X_15288_ _15284_/Y _15287_/Y _15284_/Y _15287_/Y VGND VGND VPWR VPWR _15289_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_125_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14239_ _14239_/A VGND VGND VPWR VPWR _14239_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08800_ _09213_/A VGND VGND VPWR VPWR _10014_/A sky130_fd_sc_hd__buf_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _10081_/A _09778_/Y _09779_/Y VGND VGND VPWR VPWR _09782_/B sky130_fd_sc_hd__o21ai_2
X_08731_ _08714_/Y _08729_/Y _08730_/X VGND VGND VPWR VPWR _08731_/Y sky130_fd_sc_hd__o21ai_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08662_ _08662_/A _08662_/B VGND VGND VPWR VPWR _09677_/A sky130_fd_sc_hd__or2_1
XFILLER_93_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08593_ _08592_/Y _08423_/X _08592_/Y _08423_/X VGND VGND VPWR VPWR _08596_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09214_ _09856_/A VGND VGND VPWR VPWR _09728_/A sky130_fd_sc_hd__inv_2
XFILLER_10_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09145_ _09145_/A VGND VGND VPWR VPWR _09145_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09076_ _10013_/B _09076_/B VGND VGND VPWR VPWR _09077_/B sky130_fd_sc_hd__or2_1
XFILLER_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09978_ _09978_/A _09978_/B VGND VGND VPWR VPWR _09978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08929_ _08929_/A _08929_/B VGND VGND VPWR VPWR _10287_/A sky130_fd_sc_hd__or2_1
XFILLER_92_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11940_ _13697_/A _11907_/B _11907_/Y VGND VGND VPWR VPWR _11940_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11871_ _13629_/A _11843_/B _11843_/Y VGND VGND VPWR VPWR _11871_/Y sky130_fd_sc_hd__o21ai_1
X_14590_ _15243_/A VGND VGND VPWR VPWR _14665_/A sky130_fd_sc_hd__buf_1
XFILLER_72_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13610_ _13610_/A VGND VGND VPWR VPWR _13610_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10822_ _12082_/A _10964_/B _10821_/Y VGND VGND VPWR VPWR _10823_/A sky130_fd_sc_hd__o21ai_2
XFILLER_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10753_ _13677_/A _10629_/B _10629_/Y VGND VGND VPWR VPWR _10753_/Y sky130_fd_sc_hd__o21ai_1
X_13541_ _15046_/A _13504_/B _13504_/Y _13540_/X VGND VGND VPWR VPWR _13541_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16260_ _16260_/A _16260_/B VGND VGND VPWR VPWR _16260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13472_ _13457_/X _13471_/X _13457_/X _13471_/X VGND VGND VPWR VPWR _14368_/A sky130_fd_sc_hd__a2bb2o_4
X_15211_ _15211_/A _15211_/B VGND VGND VPWR VPWR _15211_/Y sky130_fd_sc_hd__nand2_1
X_10684_ _11992_/A _10811_/B _10683_/Y VGND VGND VPWR VPWR _10685_/A sky130_fd_sc_hd__o21ai_2
XFILLER_9_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16191_ _15808_/X _16190_/X _15808_/X _16190_/X VGND VGND VPWR VPWR _16192_/B sky130_fd_sc_hd__a2bb2o_1
X_12423_ _12423_/A _12423_/B VGND VGND VPWR VPWR _12423_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12354_ _12303_/A _12303_/B _12303_/Y _12517_/A VGND VGND VPWR VPWR _12509_/A sky130_fd_sc_hd__a2bb2o_1
X_15142_ _15088_/X _15141_/Y _15088_/X _15141_/Y VGND VGND VPWR VPWR _15143_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15073_ _15073_/A _15034_/X VGND VGND VPWR VPWR _15073_/X sky130_fd_sc_hd__or2b_1
X_11305_ _13504_/A _11304_/B _11304_/X _11131_/X VGND VGND VPWR VPWR _11305_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14024_ _14109_/A _14024_/B VGND VGND VPWR VPWR _14024_/X sky130_fd_sc_hd__and2_1
X_12285_ _13793_/A _12362_/B _12284_/Y VGND VGND VPWR VPWR _12285_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11236_ _12227_/A _11236_/B VGND VGND VPWR VPWR _11236_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11167_ _12254_/A _11288_/B VGND VGND VPWR VPWR _11167_/Y sky130_fd_sc_hd__nand2_1
X_10118_ _10118_/A _10118_/B VGND VGND VPWR VPWR _10119_/A sky130_fd_sc_hd__or2_1
X_15975_ _14163_/X _15853_/A _14163_/X _15853_/A VGND VGND VPWR VPWR _15984_/B sky130_fd_sc_hd__a2bb2o_1
X_11098_ _11302_/A VGND VGND VPWR VPWR _12259_/A sky130_fd_sc_hd__buf_1
X_14926_ _15550_/A _14926_/B VGND VGND VPWR VPWR _14926_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10049_ _10049_/A _10079_/B VGND VGND VPWR VPWR _10049_/X sky130_fd_sc_hd__and2_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14857_ _14858_/A _14858_/B VGND VGND VPWR VPWR _14859_/A sky130_fd_sc_hd__and2_1
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14788_ _14788_/A _14735_/X VGND VGND VPWR VPWR _14788_/X sky130_fd_sc_hd__or2b_1
X_13808_ _13770_/X _13807_/X _13770_/X _13807_/X VGND VGND VPWR VPWR _13854_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13739_ _13739_/A _13693_/X VGND VGND VPWR VPWR _13739_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16458_ _08229_/A _16458_/D VGND VGND VPWR VPWR _16458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16389_ _16385_/X _16388_/Y _16385_/X _16388_/Y VGND VGND VPWR VPWR _16389_/X sky130_fd_sc_hd__a2bb2o_1
X_15409_ _15453_/A _15407_/X _15408_/X VGND VGND VPWR VPWR _15409_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09901_ _09901_/A _09900_/Y VGND VGND VPWR VPWR _09903_/B sky130_fd_sc_hd__or2b_1
XFILLER_113_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09832_ _09832_/A _09832_/B VGND VGND VPWR VPWR _09833_/A sky130_fd_sc_hd__nand2_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _09763_/A VGND VGND VPWR VPWR _09779_/A sky130_fd_sc_hd__inv_2
XFILLER_74_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _08714_/A _08714_/B VGND VGND VPWR VPWR _08714_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09694_ _08605_/X _09696_/B _08605_/X _09696_/B VGND VGND VPWR VPWR _09695_/B sky130_fd_sc_hd__a2bb2o_1
Xrebuffer10 rebuffer11/X VGND VGND VPWR VPWR rebuffer9/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_27_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer21 rebuffer22/X VGND VGND VPWR VPWR rebuffer21/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer32 _16316_/A VGND VGND VPWR VPWR _16381_/A1 sky130_fd_sc_hd__dlygate4sd1_1
X_08645_ _08645_/A VGND VGND VPWR VPWR _08645_/X sky130_fd_sc_hd__buf_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _08589_/A _08576_/B VGND VGND VPWR VPWR _09454_/B sky130_fd_sc_hd__or2_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09128_ _09424_/A _09131_/B VGND VGND VPWR VPWR _09128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09059_ _08806_/Y _09047_/A _08806_/A _09047_/Y VGND VGND VPWR VPWR _10015_/B sky130_fd_sc_hd__o22a_1
XFILLER_2_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12070_ _12068_/Y _12069_/Y _12008_/Y VGND VGND VPWR VPWR _12161_/A sky130_fd_sc_hd__o21ai_2
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11021_ _11021_/A VGND VGND VPWR VPWR _13552_/A sky130_fd_sc_hd__buf_1
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15760_ _14910_/A _14910_/B _14910_/Y VGND VGND VPWR VPWR _15760_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12972_ _12937_/X _12971_/Y _12937_/X _12971_/Y VGND VGND VPWR VPWR _13026_/B sky130_fd_sc_hd__a2bb2o_1
X_15691_ _15549_/X _15690_/X _15549_/X _15690_/X VGND VGND VPWR VPWR _15692_/B sky130_fd_sc_hd__a2bb2o_1
X_14711_ _14727_/A _14727_/B VGND VGND VPWR VPWR _14804_/A sky130_fd_sc_hd__and2_1
XFILLER_45_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11923_ _10685_/A _11922_/A _10685_/Y _11992_/B VGND VGND VPWR VPWR _11925_/B sky130_fd_sc_hd__o22a_1
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14642_ _15270_/A _14572_/B _14572_/Y VGND VGND VPWR VPWR _14642_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11854_ _11854_/A _11854_/B VGND VGND VPWR VPWR _11854_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10805_ _10079_/A _10804_/Y _09968_/Y _10804_/A _10957_/A VGND VGND VPWR VPWR _11988_/A
+ sky130_fd_sc_hd__o221a_1
X_14573_ _13096_/X _14571_/Y _14572_/Y VGND VGND VPWR VPWR _14573_/X sky130_fd_sc_hd__o21a_1
X_11785_ _11785_/A _11784_/X VGND VGND VPWR VPWR _11785_/X sky130_fd_sc_hd__or2b_1
XFILLER_41_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16312_ _16457_/X VGND VGND VPWR VPWR _16312_/Y sky130_fd_sc_hd__inv_2
X_10736_ _12990_/A _10635_/B _10635_/Y VGND VGND VPWR VPWR _10736_/Y sky130_fd_sc_hd__o21ai_1
X_13524_ _10317_/X _13483_/X _10317_/X _13483_/X VGND VGND VPWR VPWR _13525_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_40_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16243_ _16243_/A _16384_/B VGND VGND VPWR VPWR _16244_/A sky130_fd_sc_hd__or2_1
X_13455_ _14068_/A _13309_/B _13309_/Y _13373_/X VGND VGND VPWR VPWR _13455_/Y sky130_fd_sc_hd__o2bb2ai_1
X_10667_ _10077_/A _10666_/Y _09969_/Y _10666_/A _10957_/A VGND VGND VPWR VPWR _11916_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_127_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16174_ _16112_/A _15813_/B _15813_/Y VGND VGND VPWR VPWR _16174_/X sky130_fd_sc_hd__o21a_1
X_12406_ _12356_/X _12405_/Y _12356_/X _12405_/Y VGND VGND VPWR VPWR _12407_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13386_ _13366_/X _13385_/X _13366_/X _13385_/X VGND VGND VPWR VPWR _13442_/B sky130_fd_sc_hd__a2bb2o_1
X_10598_ _11839_/A _10529_/B _10529_/Y VGND VGND VPWR VPWR _10598_/Y sky130_fd_sc_hd__o21ai_1
X_15125_ _15125_/A _15125_/B VGND VGND VPWR VPWR _15125_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12337_ _12221_/A _12221_/B _12221_/Y VGND VGND VPWR VPWR _12337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15056_ _15045_/X _15055_/X _15045_/X _15055_/X VGND VGND VPWR VPWR _15057_/B sky130_fd_sc_hd__a2bb2o_1
X_12268_ _12268_/A _12268_/B VGND VGND VPWR VPWR _12268_/Y sky130_fd_sc_hd__nor2_1
X_11219_ _11219_/A _11219_/B VGND VGND VPWR VPWR _13337_/A sky130_fd_sc_hd__or2_1
X_14007_ _15418_/A _13960_/B _13960_/Y VGND VGND VPWR VPWR _14007_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12199_ _13894_/A _12200_/B VGND VGND VPWR VPWR _12201_/A sky130_fd_sc_hd__and2_1
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15958_ _15958_/A _15958_/B VGND VGND VPWR VPWR _15958_/X sky130_fd_sc_hd__or2_1
XFILLER_83_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14909_ _14898_/Y _14907_/X _14908_/Y VGND VGND VPWR VPWR _14909_/X sky130_fd_sc_hd__o21a_1
X_15889_ _15880_/Y _15887_/X _15888_/Y VGND VGND VPWR VPWR _15889_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08430_ _08429_/A _08333_/Y _08429_/Y _08333_/A _08441_/A VGND VGND VPWR VPWR _09209_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_91_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08361_ _08361_/A VGND VGND VPWR VPWR _08361_/Y sky130_fd_sc_hd__inv_2
X_08292_ _08321_/A input19/X _08322_/A _08324_/A VGND VGND VPWR VPWR _08319_/A sky130_fd_sc_hd__o22a_1
XFILLER_32_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09815_ _09810_/X _08830_/A _09810_/X _08830_/A VGND VGND VPWR VPWR _09819_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09746_ _09348_/B _09743_/X _08512_/X VGND VGND VPWR VPWR _09791_/B sky130_fd_sc_hd__o21a_1
XFILLER_27_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09677_/A _09677_/B VGND VGND VPWR VPWR _09681_/B sky130_fd_sc_hd__and2_1
XFILLER_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08628_ _08634_/A VGND VGND VPWR VPWR _09458_/B sky130_fd_sc_hd__buf_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08559_ _08558_/A _08439_/Y _08558_/Y _08439_/A VGND VGND VPWR VPWR _10117_/B sky130_fd_sc_hd__o22a_1
X_11570_ _14149_/A VGND VGND VPWR VPWR _12494_/A sky130_fd_sc_hd__inv_2
XFILLER_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10521_ _10521_/A _10622_/C VGND VGND VPWR VPWR _10522_/A sky130_fd_sc_hd__or2_1
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13240_ _14735_/A _13291_/B VGND VGND VPWR VPWR _13240_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10452_ _10449_/Y _12698_/A _10368_/X _10451_/Y VGND VGND VPWR VPWR _10452_/X sky130_fd_sc_hd__o22a_1
X_13171_ _13188_/A _13188_/B VGND VGND VPWR VPWR _13171_/Y sky130_fd_sc_hd__nor2_1
X_10383_ _10252_/A _10252_/B _10252_/Y VGND VGND VPWR VPWR _10384_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12122_ _13918_/A _12143_/B VGND VGND VPWR VPWR _12219_/A sky130_fd_sc_hd__and2_1
XFILLER_2_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12053_ _12053_/A _12053_/B VGND VGND VPWR VPWR _12053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11004_ _11004_/A _11003_/X VGND VGND VPWR VPWR _11004_/X sky130_fd_sc_hd__or2b_1
XFILLER_77_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15812_ _15743_/Y _15810_/X _15811_/Y VGND VGND VPWR VPWR _15812_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15743_ _16110_/A _15811_/B VGND VGND VPWR VPWR _15743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12955_ _14944_/A _12947_/B _12947_/Y VGND VGND VPWR VPWR _12955_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11906_ _11906_/A VGND VGND VPWR VPWR _11906_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15674_ _15630_/Y _15672_/X _15673_/Y VGND VGND VPWR VPWR _15674_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12886_ _12849_/X _12885_/Y _12849_/X _12885_/Y VGND VGND VPWR VPWR _12936_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _14581_/X _14624_/Y _14581_/X _14624_/Y VGND VGND VPWR VPWR _14654_/B sky130_fd_sc_hd__a2bb2o_1
X_11837_ _11837_/A _11837_/B VGND VGND VPWR VPWR _11837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _15261_/A VGND VGND VPWR VPWR _14578_/A sky130_fd_sc_hd__buf_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11768_ _12769_/A _11799_/A _11767_/Y VGND VGND VPWR VPWR _11768_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10719_ _10640_/A _10718_/Y _10640_/A _10718_/Y VGND VGND VPWR VPWR _10720_/B sky130_fd_sc_hd__a2bb2o_1
X_13507_ _13507_/A _13507_/B VGND VGND VPWR VPWR _13507_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14487_ _14466_/X _14486_/Y _14466_/X _14486_/Y VGND VGND VPWR VPWR _14518_/B sky130_fd_sc_hd__a2bb2o_1
X_11699_ _13979_/A VGND VGND VPWR VPWR _15556_/A sky130_fd_sc_hd__buf_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16226_ _16094_/A _15794_/B _15794_/Y VGND VGND VPWR VPWR _16228_/A sky130_fd_sc_hd__o21ai_1
X_13438_ _13438_/A _13438_/B VGND VGND VPWR VPWR _13438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer1 rebuffer2/X VGND VGND VPWR VPWR _11606_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_127_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16157_ _16388_/A _16157_/B VGND VGND VPWR VPWR _16268_/A sky130_fd_sc_hd__or2_1
XFILLER_115_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13369_ _13369_/A _13369_/B VGND VGND VPWR VPWR _13369_/X sky130_fd_sc_hd__or2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16088_ _16029_/X _16087_/Y _16029_/X _16087_/Y VGND VGND VPWR VPWR _16223_/A sky130_fd_sc_hd__a2bb2o_1
X_15108_ _15107_/A _15107_/B _15107_/Y VGND VGND VPWR VPWR _15108_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15039_ _15067_/A _15037_/X _15038_/X VGND VGND VPWR VPWR _15039_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09600_ _09983_/A VGND VGND VPWR VPWR _09984_/A sky130_fd_sc_hd__buf_1
XFILLER_49_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09531_ _09531_/A _09531_/B VGND VGND VPWR VPWR _09532_/A sky130_fd_sc_hd__or2_1
XFILLER_64_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09462_ _10018_/A _09462_/B VGND VGND VPWR VPWR _09462_/X sky130_fd_sc_hd__or2_1
XFILLER_52_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09393_ _09393_/A VGND VGND VPWR VPWR _09393_/X sky130_fd_sc_hd__clkbuf_2
X_08413_ _09225_/B _08408_/Y _09252_/A VGND VGND VPWR VPWR _08413_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08344_ _08344_/A VGND VGND VPWR VPWR _08344_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08275_ _08275_/A input10/X VGND VGND VPWR VPWR _08387_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09729_ _08580_/X _09731_/B _08580_/X _09731_/B VGND VGND VPWR VPWR _09730_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12740_ _12714_/X _12739_/X _12714_/X _12739_/X VGND VGND VPWR VPWR _12775_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12671_ _11140_/Y _12670_/Y _10976_/Y VGND VGND VPWR VPWR _12672_/A sky130_fd_sc_hd__o21ai_1
X_15390_ _15331_/A _15331_/B _15331_/Y VGND VGND VPWR VPWR _15390_/Y sky130_fd_sc_hd__o21ai_1
X_14410_ _14410_/A VGND VGND VPWR VPWR _15347_/A sky130_fd_sc_hd__buf_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11622_ _11617_/Y _11621_/Y _11617_/Y _11621_/Y VGND VGND VPWR VPWR _11623_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14341_ _14353_/A _14341_/B VGND VGND VPWR VPWR _15954_/A sky130_fd_sc_hd__or2_1
XFILLER_128_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11553_ _12397_/A VGND VGND VPWR VPWR _14832_/A sky130_fd_sc_hd__buf_1
XFILLER_7_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14272_ _15860_/A _14272_/B VGND VGND VPWR VPWR _14272_/Y sky130_fd_sc_hd__nand2_1
X_10504_ _10405_/A _10409_/B _10405_/A _10409_/B VGND VGND VPWR VPWR _10504_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11484_ _11583_/A _11484_/B VGND VGND VPWR VPWR _13206_/A sky130_fd_sc_hd__or2_2
X_16011_ _16011_/A _15956_/X VGND VGND VPWR VPWR _16011_/X sky130_fd_sc_hd__or2b_1
X_13223_ _13202_/A _13202_/B _13202_/Y VGND VGND VPWR VPWR _13223_/Y sky130_fd_sc_hd__o21ai_1
X_10435_ _13564_/A _10400_/B _10400_/X _10434_/X VGND VGND VPWR VPWR _10435_/X sky130_fd_sc_hd__o22a_1
XFILLER_124_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13154_ _15246_/A _13117_/B _13117_/Y VGND VGND VPWR VPWR _13154_/Y sky130_fd_sc_hd__o21ai_1
X_12105_ _13200_/A _12155_/B _12104_/Y VGND VGND VPWR VPWR _12105_/Y sky130_fd_sc_hd__o21ai_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10366_ _11757_/A VGND VGND VPWR VPWR _11750_/A sky130_fd_sc_hd__inv_2
XFILLER_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13085_ _13085_/A _13016_/X VGND VGND VPWR VPWR _13085_/X sky130_fd_sc_hd__or2b_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _10325_/B VGND VGND VPWR VPWR _12701_/A sky130_fd_sc_hd__inv_2
X_12036_ _11965_/X _12035_/Y _11965_/X _12035_/Y VGND VGND VPWR VPWR _12051_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13987_ _13862_/X _13884_/A _13883_/X VGND VGND VPWR VPWR _13987_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15726_ _15546_/A _14922_/B _14922_/Y VGND VGND VPWR VPWR _15726_/X sky130_fd_sc_hd__o21a_1
X_12938_ _12938_/A _12938_/B VGND VGND VPWR VPWR _12938_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15657_ _15509_/A _15509_/B _15510_/A VGND VGND VPWR VPWR _15658_/A sky130_fd_sc_hd__o21ai_1
XFILLER_61_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14608_ _14665_/A _14665_/B _14607_/Y VGND VGND VPWR VPWR _14608_/Y sky130_fd_sc_hd__o21ai_1
X_12869_ _12858_/A _12858_/B _12858_/Y VGND VGND VPWR VPWR _12869_/Y sky130_fd_sc_hd__o21ai_1
X_15588_ _15700_/A _15588_/B VGND VGND VPWR VPWR _16046_/A sky130_fd_sc_hd__or2_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14539_ _14588_/A _14588_/B VGND VGND VPWR VPWR _14539_/Y sky130_fd_sc_hd__nor2_1
X_16209_ _16207_/A _16208_/A _16207_/Y _16208_/Y _15832_/A VGND VGND VPWR VPWR _16255_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08962_ _10017_/A VGND VGND VPWR VPWR _08962_/X sky130_fd_sc_hd__buf_1
XFILLER_69_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08893_ _10013_/A VGND VGND VPWR VPWR _08893_/X sky130_fd_sc_hd__buf_1
XFILLER_111_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09514_ _09488_/A _09488_/B _09488_/Y _09513_/X VGND VGND VPWR VPWR _09514_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09445_ _09445_/A VGND VGND VPWR VPWR _10926_/A sky130_fd_sc_hd__clkbuf_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09376_ _10239_/A VGND VGND VPWR VPWR _09377_/B sky130_fd_sc_hd__buf_1
X_08327_ _08327_/A _08327_/B VGND VGND VPWR VPWR _08328_/A sky130_fd_sc_hd__or2_1
XFILLER_20_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08258_ input15/X VGND VGND VPWR VPWR _08336_/A sky130_fd_sc_hd__inv_2
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10220_ _11745_/A VGND VGND VPWR VPWR _10224_/A sky130_fd_sc_hd__inv_2
XFILLER_106_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10151_ _10151_/A _10151_/B VGND VGND VPWR VPWR _10151_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10082_ _10046_/X _10080_/X _10967_/B VGND VGND VPWR VPWR _10082_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13910_ _13910_/A VGND VGND VPWR VPWR _15408_/A sky130_fd_sc_hd__buf_1
XFILLER_87_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14890_ _14802_/A _14802_/B _14802_/A _14802_/B VGND VGND VPWR VPWR _14890_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13841_ _13832_/Y _13839_/X _13840_/Y VGND VGND VPWR VPWR _13841_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13772_ _13807_/A _13770_/X _13771_/X VGND VGND VPWR VPWR _13772_/X sky130_fd_sc_hd__o21a_1
X_10984_ _12172_/A VGND VGND VPWR VPWR _12688_/A sky130_fd_sc_hd__buf_1
XFILLER_28_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15511_ _15509_/A _15509_/B _12609_/A _15510_/Y VGND VGND VPWR VPWR _15512_/B sky130_fd_sc_hd__o22a_1
X_12723_ _13458_/A _13458_/B _12722_/Y VGND VGND VPWR VPWR _12723_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15442_ _15415_/X _15441_/X _15415_/X _15441_/X VGND VGND VPWR VPWR _15443_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12654_ _13979_/A VGND VGND VPWR VPWR _14948_/A sky130_fd_sc_hd__inv_2
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12585_ _12585_/A VGND VGND VPWR VPWR _12585_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15373_ _15342_/X _15372_/X _15342_/X _15372_/X VGND VGND VPWR VPWR _15410_/B sky130_fd_sc_hd__a2bb2o_1
X_11605_ _12423_/A VGND VGND VPWR VPWR _11609_/A sky130_fd_sc_hd__inv_2
XFILLER_30_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14324_ _15960_/A _14390_/B VGND VGND VPWR VPWR _15605_/A sky130_fd_sc_hd__and2_1
X_11536_ _11620_/A _12416_/A _11535_/Y VGND VGND VPWR VPWR _11536_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14255_ _14228_/Y _14253_/Y _14254_/Y VGND VGND VPWR VPWR _14256_/A sky130_fd_sc_hd__o21ai_1
XFILLER_116_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13206_ _13206_/A _13206_/B VGND VGND VPWR VPWR _13206_/Y sky130_fd_sc_hd__nand2_1
X_11467_ _09430_/A _09185_/B _09185_/Y VGND VGND VPWR VPWR _11468_/A sky130_fd_sc_hd__o21ai_1
X_14186_ _15857_/A _14275_/B VGND VGND VPWR VPWR _14186_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10418_ _12831_/A _10355_/B _10356_/A VGND VGND VPWR VPWR _10418_/Y sky130_fd_sc_hd__o21ai_1
X_11398_ _08960_/A _08960_/B _08960_/Y VGND VGND VPWR VPWR _11399_/A sky130_fd_sc_hd__o21ai_1
XFILLER_98_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13137_ _14976_/A _13127_/B _13127_/Y VGND VGND VPWR VPWR _13137_/Y sky130_fd_sc_hd__o21ai_1
X_10349_ _10349_/A VGND VGND VPWR VPWR _10350_/B sky130_fd_sc_hd__inv_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13068_ _13068_/A VGND VGND VPWR VPWR _13767_/A sky130_fd_sc_hd__inv_2
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _12059_/A VGND VGND VPWR VPWR _13194_/A sky130_fd_sc_hd__buf_1
XFILLER_93_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15709_ _15728_/A _15709_/B VGND VGND VPWR VPWR _16123_/A sky130_fd_sc_hd__or2_1
XFILLER_81_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09230_ _09230_/A _09800_/A VGND VGND VPWR VPWR _09230_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09161_ _08708_/Y _09160_/Y _08746_/X VGND VGND VPWR VPWR _09161_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09092_ _09703_/A VGND VGND VPWR VPWR _09418_/A sky130_fd_sc_hd__buf_1
XFILLER_119_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09994_ _09966_/Y _09992_/Y _09993_/Y VGND VGND VPWR VPWR _11307_/A sky130_fd_sc_hd__o21ai_1
XFILLER_103_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08945_ _08844_/A _08842_/Y _08944_/X VGND VGND VPWR VPWR _08946_/A sky130_fd_sc_hd__o21ai_1
XFILLER_57_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08876_ _08876_/A _08876_/B VGND VGND VPWR VPWR _08876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09428_ _09428_/A VGND VGND VPWR VPWR _09428_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09359_ _09478_/B _09863_/A _09347_/Y _09358_/X VGND VGND VPWR VPWR _09359_/X sky130_fd_sc_hd__o22a_1
X_12370_ _12370_/A VGND VGND VPWR VPWR _12370_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11321_ _11321_/A VGND VGND VPWR VPWR _11321_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14040_ _14043_/A VGND VGND VPWR VPWR _14812_/A sky130_fd_sc_hd__buf_1
X_11252_ _13349_/A _11242_/B _11242_/Y _11251_/X VGND VGND VPWR VPWR _11252_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11183_ _13367_/A VGND VGND VPWR VPWR _14015_/A sky130_fd_sc_hd__inv_2
XFILLER_69_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10203_ _10215_/A _11243_/A VGND VGND VPWR VPWR _10282_/A sky130_fd_sc_hd__or2_2
XFILLER_106_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10134_ _10134_/A _10134_/B VGND VGND VPWR VPWR _10134_/X sky130_fd_sc_hd__or2_1
X_15991_ _15991_/A _15991_/B VGND VGND VPWR VPWR _15991_/X sky130_fd_sc_hd__or2_1
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14942_ _15171_/A _14980_/B VGND VGND VPWR VPWR _14942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10065_ _10065_/A _10065_/B VGND VGND VPWR VPWR _10065_/Y sky130_fd_sc_hd__nor2_1
X_14873_ _14782_/A _14782_/B _14782_/A _14782_/B VGND VGND VPWR VPWR _14873_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13824_ _14631_/A _13844_/B VGND VGND VPWR VPWR _13824_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13755_ _13755_/A VGND VGND VPWR VPWR _13755_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10967_ _10046_/X _10967_/B VGND VGND VPWR VPWR _10967_/X sky130_fd_sc_hd__and2b_1
X_16474_ _16474_/D _16454_/Y VGND VGND VPWR VPWR _16474_/Q sky130_fd_sc_hd__dlxtn_1
X_10898_ _13829_/A _10909_/B VGND VGND VPWR VPWR _10898_/Y sky130_fd_sc_hd__nor2_1
X_13686_ _13686_/A VGND VGND VPWR VPWR _13686_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12706_ _12706_/A _12706_/B VGND VGND VPWR VPWR _12706_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12637_ _12637_/A _12637_/B VGND VGND VPWR VPWR _12637_/X sky130_fd_sc_hd__or2_1
X_15425_ _15425_/A _15425_/B VGND VGND VPWR VPWR _15425_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12568_ _12564_/Y _12567_/Y _12564_/A _12567_/A _11706_/A VGND VGND VPWR VPWR _12623_/A
+ sky130_fd_sc_hd__o221a_1
X_15356_ _15422_/A _15422_/B VGND VGND VPWR VPWR _15356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12499_ _12499_/A VGND VGND VPWR VPWR _12500_/A sky130_fd_sc_hd__clkbuf_2
X_14307_ _13442_/A _13442_/B _13442_/Y VGND VGND VPWR VPWR _14307_/X sky130_fd_sc_hd__o21a_1
X_15287_ _15287_/A _15287_/B VGND VGND VPWR VPWR _15287_/Y sky130_fd_sc_hd__nor2_1
X_11519_ _11518_/Y _11315_/X _11324_/Y VGND VGND VPWR VPWR _11519_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14238_ _15509_/A _14082_/B _14082_/Y VGND VGND VPWR VPWR _14239_/A sky130_fd_sc_hd__a21oi_1
X_14169_ _14140_/X _14168_/Y _14140_/X _14168_/Y VGND VGND VPWR VPWR _14170_/B sky130_fd_sc_hd__a2bb2oi_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08730_ _09213_/A _09454_/B VGND VGND VPWR VPWR _08730_/X sky130_fd_sc_hd__or2_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08661_ _08919_/A VGND VGND VPWR VPWR _09235_/A sky130_fd_sc_hd__buf_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08592_ _08592_/A VGND VGND VPWR VPWR _08592_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09213_ _09213_/A _09213_/B VGND VGND VPWR VPWR _09856_/A sky130_fd_sc_hd__or2_2
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09144_ _09432_/A _09175_/B _09143_/Y VGND VGND VPWR VPWR _09145_/A sky130_fd_sc_hd__o21ai_1
XFILLER_108_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09075_ _10014_/B _09075_/B VGND VGND VPWR VPWR _09076_/B sky130_fd_sc_hd__or2_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09977_ _09977_/A _09978_/B VGND VGND VPWR VPWR _09977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08928_ _08928_/A VGND VGND VPWR VPWR _08929_/B sky130_fd_sc_hd__inv_2
XFILLER_72_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08859_ _09500_/A _08834_/A _08836_/Y _08955_/A VGND VGND VPWR VPWR _08859_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11870_ _11907_/A _11907_/B VGND VGND VPWR VPWR _11870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10821_ _12082_/A _10964_/B VGND VGND VPWR VPWR _10821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10752_ _11892_/A VGND VGND VPWR VPWR _13677_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13540_ _15044_/A _13507_/B _13507_/Y _13539_/X VGND VGND VPWR VPWR _13540_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13471_ _13459_/X _13470_/X _13459_/X _13470_/X VGND VGND VPWR VPWR _13471_/X sky130_fd_sc_hd__a2bb2o_2
X_15210_ _15147_/X _15209_/Y _15147_/X _15209_/Y VGND VGND VPWR VPWR _15211_/B sky130_fd_sc_hd__a2bb2o_1
X_12422_ _12422_/A VGND VGND VPWR VPWR _12422_/Y sky130_fd_sc_hd__inv_2
X_10683_ _11992_/A _10811_/B VGND VGND VPWR VPWR _10683_/Y sky130_fd_sc_hd__nand2_1
X_16190_ _16108_/A _15809_/B _15809_/Y VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__o21a_1
X_12353_ _12306_/A _12306_/B _12306_/Y _12525_/A VGND VGND VPWR VPWR _12517_/A sky130_fd_sc_hd__a2bb2o_1
X_15141_ _15084_/A _15084_/B _15084_/Y VGND VGND VPWR VPWR _15141_/Y sky130_fd_sc_hd__o21ai_1
X_12284_ _12362_/A _12362_/B VGND VGND VPWR VPWR _12284_/Y sky130_fd_sc_hd__nand2_1
X_15072_ _15072_/A _15072_/B VGND VGND VPWR VPWR _15072_/Y sky130_fd_sc_hd__nand2_1
X_11304_ _12170_/A _11304_/B VGND VGND VPWR VPWR _11304_/X sky130_fd_sc_hd__and2_1
XFILLER_5_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14023_ _13949_/X _14022_/Y _13949_/X _14022_/Y VGND VGND VPWR VPWR _14024_/B sky130_fd_sc_hd__a2bb2o_1
X_11235_ _11077_/X _11234_/X _11077_/X _11234_/X VGND VGND VPWR VPWR _11236_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11166_ _11123_/X _11165_/Y _11123_/X _11165_/Y VGND VGND VPWR VPWR _11288_/B sky130_fd_sc_hd__a2bb2o_1
X_15974_ _15974_/A VGND VGND VPWR VPWR _15984_/A sky130_fd_sc_hd__inv_2
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10117_ _10117_/A _10117_/B VGND VGND VPWR VPWR _10118_/A sky130_fd_sc_hd__or2_1
X_11097_ _11096_/A _11096_/B _11096_/Y _09393_/X VGND VGND VPWR VPWR _11302_/A sky130_fd_sc_hd__o211a_1
X_14925_ _14871_/Y _14923_/X _14924_/Y VGND VGND VPWR VPWR _14925_/X sky130_fd_sc_hd__o21a_1
X_10048_ _10025_/X _10047_/Y _10025_/X _10047_/Y VGND VGND VPWR VPWR _10079_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14856_ _14831_/X _14855_/Y _14831_/X _14855_/Y VGND VGND VPWR VPWR _14858_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08231__1 _16357_/A VGND VGND VPWR VPWR _16358_/A sky130_fd_sc_hd__inv_2
X_14787_ _15452_/A VGND VGND VPWR VPWR _14790_/A sky130_fd_sc_hd__buf_1
X_13807_ _13807_/A _13771_/X VGND VGND VPWR VPWR _13807_/X sky130_fd_sc_hd__or2b_1
XFILLER_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13738_ _13765_/A _13765_/B VGND VGND VPWR VPWR _13816_/A sky130_fd_sc_hd__and2_1
X_11999_ _12080_/B _11998_/X _12080_/B _11998_/X VGND VGND VPWR VPWR _12076_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16457_ _16395_/A _16248_/B _16457_/S VGND VGND VPWR VPWR _16457_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13669_ _13624_/A _13668_/Y _13624_/A _13668_/Y VGND VGND VPWR VPWR _13693_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16388_ _16388_/A _16388_/B VGND VGND VPWR VPWR _16388_/Y sky130_fd_sc_hd__nor2_1
X_15408_ _15408_/A _15408_/B VGND VGND VPWR VPWR _15408_/X sky130_fd_sc_hd__or2_1
X_15339_ _15339_/A _15339_/B VGND VGND VPWR VPWR _15339_/X sky130_fd_sc_hd__or2_1
X_09900_ _09898_/A _09898_/B _09899_/Y VGND VGND VPWR VPWR _09900_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _09829_/A _09829_/B _09830_/Y _08931_/Y VGND VGND VPWR VPWR _09832_/B sky130_fd_sc_hd__o22a_1
XFILLER_112_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _10046_/A VGND VGND VPWR VPWR _10081_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08713_/A _08713_/B VGND VGND VPWR VPWR _08713_/X sky130_fd_sc_hd__or2_1
XFILLER_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09693_ _09693_/A _09693_/B VGND VGND VPWR VPWR _09696_/B sky130_fd_sc_hd__or2_1
Xrebuffer11 rebuffer12/X VGND VGND VPWR VPWR rebuffer11/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_82_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer33 _08358_/A VGND VGND VPWR VPWR _08393_/A1 sky130_fd_sc_hd__dlygate4sd1_1
X_08644_ _09458_/A _09228_/B _09228_/A _08386_/Y VGND VGND VPWR VPWR _08645_/A sky130_fd_sc_hd__o22a_1
Xrebuffer22 rebuffer23/X VGND VGND VPWR VPWR rebuffer22/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08575_ _08574_/A _08338_/Y _08574_/Y _08338_/A VGND VGND VPWR VPWR _08576_/B sky130_fd_sc_hd__o22a_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09127_ _09088_/Y _09125_/Y _09126_/Y VGND VGND VPWR VPWR _09131_/B sky130_fd_sc_hd__o21ai_1
XFILLER_108_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09058_ _08798_/X _09048_/Y _08798_/X _09048_/Y VGND VGND VPWR VPWR _10014_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11020_ _13906_/A _11089_/B VGND VGND VPWR VPWR _11204_/A sky130_fd_sc_hd__and2_1
XFILLER_2_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12971_ _14532_/A _12938_/B _12938_/Y VGND VGND VPWR VPWR _12971_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15690_ _15494_/X _15690_/B VGND VGND VPWR VPWR _15690_/X sky130_fd_sc_hd__and2b_1
X_14710_ _14649_/X _14709_/Y _14649_/X _14709_/Y VGND VGND VPWR VPWR _14727_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11922_ _11922_/A VGND VGND VPWR VPWR _11992_/B sky130_fd_sc_hd__inv_2
X_14641_ _14646_/A _14646_/B VGND VGND VPWR VPWR _14716_/A sky130_fd_sc_hd__and2_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11853_ _11852_/A _11852_/B _11852_/X _11810_/B VGND VGND VPWR VPWR _11918_/B sky130_fd_sc_hd__a22o_1
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10804_ _10804_/A VGND VGND VPWR VPWR _10804_/Y sky130_fd_sc_hd__inv_2
X_16311_ _16318_/A _16318_/B VGND VGND VPWR VPWR _16311_/Y sky130_fd_sc_hd__nor2_1
X_14572_ _15270_/A _14572_/B VGND VGND VPWR VPWR _14572_/Y sky130_fd_sc_hd__nand2_1
X_11784_ _13530_/A _11784_/B VGND VGND VPWR VPWR _11784_/X sky130_fd_sc_hd__or2_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10735_ _10735_/A VGND VGND VPWR VPWR _12990_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13523_ _13525_/A VGND VGND VPWR VPWR _15032_/A sky130_fd_sc_hd__buf_1
XFILLER_9_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16242_ _15781_/A _15781_/B _16241_/Y VGND VGND VPWR VPWR _16384_/B sky130_fd_sc_hd__a21oi_1
XFILLER_127_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13454_ _13451_/X _13453_/Y _13451_/X _13453_/Y VGND VGND VPWR VPWR _13454_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10666_ _10666_/A VGND VGND VPWR VPWR _10666_/Y sky130_fd_sc_hd__inv_2
X_16173_ _16189_/A _16173_/B VGND VGND VPWR VPWR _16264_/A sky130_fd_sc_hd__or2_1
XFILLER_126_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12405_ _12404_/A _12404_/B _12404_/Y VGND VGND VPWR VPWR _12405_/Y sky130_fd_sc_hd__o21ai_1
X_13385_ _13385_/A _13367_/X VGND VGND VPWR VPWR _13385_/X sky130_fd_sc_hd__or2b_1
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15124_ _15094_/X _15123_/Y _15094_/X _15123_/Y VGND VGND VPWR VPWR _15125_/B sky130_fd_sc_hd__a2bb2o_1
X_10597_ _09963_/Y _10596_/A _09963_/A _10596_/Y _09797_/A VGND VGND VPWR VPWR _10735_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12336_ _13396_/A _12339_/B VGND VGND VPWR VPWR _12336_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15055_ _15055_/A _15046_/X VGND VGND VPWR VPWR _15055_/X sky130_fd_sc_hd__or2b_1
X_12267_ _12686_/A _12266_/B _12266_/X _12179_/B VGND VGND VPWR VPWR _12373_/B sky130_fd_sc_hd__a22o_1
X_11218_ _12218_/A _11218_/B VGND VGND VPWR VPWR _11218_/Y sky130_fd_sc_hd__nand2_1
X_14006_ _14066_/A _14066_/B VGND VGND VPWR VPWR _14141_/A sky130_fd_sc_hd__and2_1
X_12198_ _12156_/X _12197_/Y _12156_/X _12197_/Y VGND VGND VPWR VPWR _12200_/B sky130_fd_sc_hd__a2bb2o_1
X_11149_ _11148_/A _11147_/Y _11148_/Y _11147_/A _11526_/A VGND VGND VPWR VPWR _11314_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_110_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15957_ _16011_/A _15955_/X _15956_/X VGND VGND VPWR VPWR _15957_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15888_ _15888_/A _15888_/B VGND VGND VPWR VPWR _15888_/Y sky130_fd_sc_hd__nand2_1
X_14908_ _14908_/A _14908_/B VGND VGND VPWR VPWR _14908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14839_ _15051_/A _12370_/Y _12276_/Y _14752_/X VGND VGND VPWR VPWR _14839_/X sky130_fd_sc_hd__o22a_1
XFILLER_24_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08360_ input9/X _08279_/B _08359_/X VGND VGND VPWR VPWR _08361_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08291_ _08326_/A input33/X _08327_/A _08329_/A VGND VGND VPWR VPWR _08324_/A sky130_fd_sc_hd__o22a_1
XFILLER_118_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09814_ _09811_/X _08822_/A _09811_/X _08822_/A VGND VGND VPWR VPWR _09820_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09745_ _09745_/A _09745_/B VGND VGND VPWR VPWR _09791_/A sky130_fd_sc_hd__or2_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _11939_/A VGND VGND VPWR VPWR _13063_/A sky130_fd_sc_hd__buf_1
XFILLER_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08627_ _08650_/A _08627_/B VGND VGND VPWR VPWR _08634_/A sky130_fd_sc_hd__or2_1
XFILLER_82_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08558_ _08558_/A VGND VGND VPWR VPWR _08558_/Y sky130_fd_sc_hd__inv_2
X_08489_ _08336_/A _08260_/B _08475_/Y _08574_/A VGND VGND VPWR VPWR _08561_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10520_ _10903_/A _11592_/A VGND VGND VPWR VPWR _10622_/C sky130_fd_sc_hd__or2_1
XFILLER_109_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10451_ _10451_/A _11764_/A VGND VGND VPWR VPWR _10451_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13170_ _13106_/X _13169_/Y _13106_/X _13169_/Y VGND VGND VPWR VPWR _13188_/B sky130_fd_sc_hd__a2bb2o_1
X_10382_ _10370_/X _10381_/Y _10370_/X _10381_/Y VGND VGND VPWR VPWR _10451_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12121_ _12054_/X _12120_/Y _12054_/X _12120_/Y VGND VGND VPWR VPWR _12143_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12052_ _12037_/Y _12050_/X _12051_/Y VGND VGND VPWR VPWR _12052_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11003_ _14410_/A _11003_/B VGND VGND VPWR VPWR _11003_/X sky130_fd_sc_hd__or2_1
XFILLER_77_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15811_ _16110_/A _15811_/B VGND VGND VPWR VPWR _15811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15742_ _15678_/X _15741_/Y _15678_/X _15741_/Y VGND VGND VPWR VPWR _15811_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12954_ _13879_/A VGND VGND VPWR VPWR _14836_/A sky130_fd_sc_hd__buf_1
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11905_ _11873_/Y _11903_/Y _11904_/Y VGND VGND VPWR VPWR _11906_/A sky130_fd_sc_hd__o21ai_1
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15673_ _15673_/A _15673_/B VGND VGND VPWR VPWR _15673_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12885_ _12850_/A _12850_/B _12850_/Y VGND VGND VPWR VPWR _12885_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14582_/A _14582_/B _14582_/Y VGND VGND VPWR VPWR _14624_/Y sky130_fd_sc_hd__o21ai_1
X_11836_ _11830_/Y _11834_/X _11835_/Y VGND VGND VPWR VPWR _11836_/X sky130_fd_sc_hd__o21a_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _14580_/A _14580_/B VGND VGND VPWR VPWR _14555_/Y sky130_fd_sc_hd__nor2_1
X_11767_ _12769_/A _11799_/A VGND VGND VPWR VPWR _11767_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10718_ _13695_/A _10641_/B _10641_/Y VGND VGND VPWR VPWR _10718_/Y sky130_fd_sc_hd__o21ai_1
X_13506_ _10986_/X _13489_/X _10986_/X _13489_/X VGND VGND VPWR VPWR _13507_/B sky130_fd_sc_hd__o2bb2a_1
X_16225_ _16223_/A _16224_/A _16223_/Y _16224_/Y _16205_/A VGND VGND VPWR VPWR _16251_/A
+ sky130_fd_sc_hd__a221o_1
X_14486_ _14467_/A _14467_/B _14467_/Y VGND VGND VPWR VPWR _14486_/Y sky130_fd_sc_hd__o21ai_1
X_11698_ _12452_/A VGND VGND VPWR VPWR _13979_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13437_ _13433_/Y _13435_/Y _13436_/Y VGND VGND VPWR VPWR _13437_/X sky130_fd_sc_hd__o21a_1
X_10649_ _11978_/A VGND VGND VPWR VPWR _13699_/A sky130_fd_sc_hd__buf_1
Xrebuffer2 rebuffer5/X VGND VGND VPWR VPWR rebuffer2/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_127_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16156_ _16113_/X _16155_/X _16113_/X _16155_/X VGND VGND VPWR VPWR _16157_/B sky130_fd_sc_hd__a2bb2oi_1
X_13368_ _13385_/A _13366_/X _13367_/X VGND VGND VPWR VPWR _13368_/X sky130_fd_sc_hd__o21a_1
X_16087_ _16030_/A _16030_/B _16030_/Y VGND VGND VPWR VPWR _16087_/Y sky130_fd_sc_hd__o21ai_1
X_12319_ _12319_/A VGND VGND VPWR VPWR _12319_/Y sky130_fd_sc_hd__inv_2
X_15107_ _15107_/A _15107_/B VGND VGND VPWR VPWR _15107_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13299_ _13299_/A VGND VGND VPWR VPWR _13299_/Y sky130_fd_sc_hd__inv_2
X_15038_ _15038_/A _15038_/B VGND VGND VPWR VPWR _15038_/X sky130_fd_sc_hd__or2_1
XFILLER_96_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09530_ _09530_/A VGND VGND VPWR VPWR _09530_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09461_ _09459_/A _08639_/B _09459_/Y _09460_/Y VGND VGND VPWR VPWR _09461_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09392_ _09392_/A VGND VGND VPWR VPWR _09393_/A sky130_fd_sc_hd__clkbuf_2
X_08412_ _08717_/A VGND VGND VPWR VPWR _09252_/A sky130_fd_sc_hd__buf_1
XFILLER_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08343_ _08343_/A VGND VGND VPWR VPWR _08343_/Y sky130_fd_sc_hd__inv_2
X_08274_ input26/X VGND VGND VPWR VPWR _08275_/A sky130_fd_sc_hd__inv_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09728_ _09728_/A _09728_/B VGND VGND VPWR VPWR _09731_/B sky130_fd_sc_hd__or2_1
XFILLER_28_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09659_ _09597_/Y _09657_/X _09658_/Y VGND VGND VPWR VPWR _09659_/X sky130_fd_sc_hd__o21a_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12670_ _12670_/A VGND VGND VPWR VPWR _12670_/Y sky130_fd_sc_hd__inv_2
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11618_/Y _12416_/A _11517_/X _11620_/Y VGND VGND VPWR VPWR _11621_/Y sky130_fd_sc_hd__o22ai_2
X_14340_ _13425_/Y _14339_/X _13425_/Y _14339_/X VGND VGND VPWR VPWR _14341_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11552_ _12397_/A _11554_/B VGND VGND VPWR VPWR _11555_/A sky130_fd_sc_hd__and2_1
X_14271_ _14271_/A VGND VGND VPWR VPWR _14271_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10503_ _11837_/A VGND VGND VPWR VPWR _13606_/A sky130_fd_sc_hd__buf_1
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11483_ _09439_/X _11482_/X _09439_/X _11482_/X VGND VGND VPWR VPWR _11484_/B sky130_fd_sc_hd__a2bb2o_1
X_16010_ _16040_/A _16040_/B VGND VGND VPWR VPWR _16010_/Y sky130_fd_sc_hd__nor2_1
X_13222_ _14674_/A VGND VGND VPWR VPWR _14741_/A sky130_fd_sc_hd__buf_1
X_10434_ _13568_/A _10409_/B _10409_/X _10433_/X VGND VGND VPWR VPWR _10434_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13153_ _13200_/A _13200_/B VGND VGND VPWR VPWR _13153_/Y sky130_fd_sc_hd__nor2_1
X_10365_ _10367_/A VGND VGND VPWR VPWR _10365_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12104_ _12104_/A _12155_/B VGND VGND VPWR VPWR _12104_/Y sky130_fd_sc_hd__nand2_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13084_ _13761_/A VGND VGND VPWR VPWR _15261_/A sky130_fd_sc_hd__buf_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10296_/A VGND VGND VPWR VPWR _10325_/A sky130_fd_sc_hd__inv_2
XFILLER_2_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12035_ _11966_/A _11966_/B _11966_/Y VGND VGND VPWR VPWR _12035_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13986_ _13986_/A _13985_/X VGND VGND VPWR VPWR _13986_/X sky130_fd_sc_hd__or2b_1
XFILLER_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15725_ _15817_/A _15817_/B VGND VGND VPWR VPWR _15725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12937_ _12887_/Y _12935_/X _12936_/Y VGND VGND VPWR VPWR _12937_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15656_ _15656_/A VGND VGND VPWR VPWR _16028_/A sky130_fd_sc_hd__inv_2
X_12868_ _12944_/A VGND VGND VPWR VPWR _14757_/A sky130_fd_sc_hd__buf_1
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14607_ _14665_/A _14665_/B VGND VGND VPWR VPWR _14607_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11819_ _11770_/A _11770_/B _11770_/A _11770_/B VGND VGND VPWR VPWR _11819_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15587_ _15545_/X _15586_/X _15545_/X _15586_/X VGND VGND VPWR VPWR _15588_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12779_/A _12779_/B _12779_/Y VGND VGND VPWR VPWR _12799_/Y sky130_fd_sc_hd__o21ai_1
X_14538_ _14523_/X _14537_/X _14523_/X _14537_/X VGND VGND VPWR VPWR _14588_/B sky130_fd_sc_hd__a2bb2o_1
X_14469_ _14469_/A _14469_/B VGND VGND VPWR VPWR _14469_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16208_ _16208_/A VGND VGND VPWR VPWR _16208_/Y sky130_fd_sc_hd__inv_2
X_16139_ _16139_/A VGND VGND VPWR VPWR _16139_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08961_ _08957_/Y _11397_/A _08960_/Y VGND VGND VPWR VPWR _08968_/A sky130_fd_sc_hd__o21ai_1
XFILLER_130_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08892_ _08686_/X _08891_/X _08686_/X _08891_/X VGND VGND VPWR VPWR _08976_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09513_ _09490_/A _09490_/B _09490_/Y _09512_/X VGND VGND VPWR VPWR _09513_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09444_ _10904_/A VGND VGND VPWR VPWR _09445_/A sky130_fd_sc_hd__clkbuf_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09375_ _09336_/X _08878_/Y _09336_/X _08878_/Y VGND VGND VPWR VPWR _10239_/A sky130_fd_sc_hd__o2bb2a_1
X_08326_ _08326_/A input33/X VGND VGND VPWR VPWR _08327_/B sky130_fd_sc_hd__nor2_1
X_08257_ input16/X _08257_/B VGND VGND VPWR VPWR _08332_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10150_ _08786_/B _10130_/B _10131_/B VGND VGND VPWR VPWR _10151_/B sky130_fd_sc_hd__a21bo_1
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10081_ _10081_/A _10081_/B VGND VGND VPWR VPWR _10967_/B sky130_fd_sc_hd__or2_1
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13840_ _14646_/A _13840_/B VGND VGND VPWR VPWR _13840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13771_ _13771_/A _13771_/B VGND VGND VPWR VPWR _13771_/X sky130_fd_sc_hd__or2_1
XFILLER_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10983_ _10981_/A _10981_/B _10981_/Y _10982_/X VGND VGND VPWR VPWR _12172_/A sky130_fd_sc_hd__o211a_1
X_15510_ _15510_/A VGND VGND VPWR VPWR _15510_/Y sky130_fd_sc_hd__inv_2
X_12722_ _13458_/A _13458_/B VGND VGND VPWR VPWR _12722_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15441_ _15441_/A _15416_/X VGND VGND VPWR VPWR _15441_/X sky130_fd_sc_hd__or2b_1
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12653_ _13985_/A VGND VGND VPWR VPWR _14976_/A sky130_fd_sc_hd__buf_1
XFILLER_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12584_ _12621_/A _12621_/B VGND VGND VPWR VPWR _14220_/A sky130_fd_sc_hd__and2_1
X_15372_ _15372_/A _15343_/X VGND VGND VPWR VPWR _15372_/X sky130_fd_sc_hd__or2b_1
X_11604_ _11604_/A _11604_/B VGND VGND VPWR VPWR _12423_/A sky130_fd_sc_hd__or2_1
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14323_ _14268_/A _14322_/Y _14268_/A _14322_/Y VGND VGND VPWR VPWR _14390_/B sky130_fd_sc_hd__a2bb2o_1
X_11535_ _11620_/A _12416_/A VGND VGND VPWR VPWR _11535_/Y sky130_fd_sc_hd__nor2_1
X_14254_ _15878_/A _14254_/B VGND VGND VPWR VPWR _14254_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11466_ _15440_/A _11353_/B _11353_/Y _11261_/X VGND VGND VPWR VPWR _11466_/X sky130_fd_sc_hd__a2bb2o_1
X_13205_ _13147_/Y _13203_/X _13204_/Y VGND VGND VPWR VPWR _13205_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14185_ _12632_/X _14184_/X _12632_/X _14184_/X VGND VGND VPWR VPWR _14275_/B sky130_fd_sc_hd__a2bb2o_1
X_10417_ _10429_/A VGND VGND VPWR VPWR _12826_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11397_ _11397_/A VGND VGND VPWR VPWR _11397_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13136_ _13139_/A VGND VGND VPWR VPWR _15289_/A sky130_fd_sc_hd__buf_1
X_10348_ _10455_/A _11711_/B VGND VGND VPWR VPWR _10349_/A sky130_fd_sc_hd__nand2_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13067_ _15249_/A _13115_/B VGND VGND VPWR VPWR _13067_/Y sky130_fd_sc_hd__nor2_1
X_10279_ _11713_/A VGND VGND VPWR VPWR _11720_/A sky130_fd_sc_hd__inv_2
XFILLER_2_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ _13196_/A _12061_/B VGND VGND VPWR VPWR _12018_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13969_ _13969_/A _13968_/X VGND VGND VPWR VPWR _13969_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15708_ _14927_/X _15707_/X _14927_/X _15707_/X VGND VGND VPWR VPWR _15709_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_74_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15639_ _15639_/A _15519_/X VGND VGND VPWR VPWR _15641_/A sky130_fd_sc_hd__or2b_1
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09160_ _09160_/A VGND VGND VPWR VPWR _09160_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09091_ _10016_/B _09073_/B _09074_/B VGND VGND VPWR VPWR _09703_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09993_ _09993_/A _09993_/B VGND VGND VPWR VPWR _09993_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08944_ _08944_/A _08944_/B VGND VGND VPWR VPWR _08944_/X sky130_fd_sc_hd__or2_1
XFILLER_88_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08875_ _08984_/A _08984_/B VGND VGND VPWR VPWR _08875_/X sky130_fd_sc_hd__and2_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09427_ _09426_/A _09433_/B _09426_/Y VGND VGND VPWR VPWR _09428_/A sky130_fd_sc_hd__o21ai_1
XFILLER_40_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09358_ _08694_/A _09862_/A _09349_/Y _09357_/X VGND VGND VPWR VPWR _09358_/X sky130_fd_sc_hd__o22a_1
X_08309_ _08309_/A VGND VGND VPWR VPWR _08309_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09289_ _09238_/A _09288_/Y _09238_/A _09288_/Y VGND VGND VPWR VPWR _10402_/A sky130_fd_sc_hd__a2bb2o_2
X_11320_ _10239_/B _10143_/B _10143_/Y VGND VGND VPWR VPWR _11321_/A sky130_fd_sc_hd__a21oi_1
XFILLER_119_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11251_ _11248_/X _11249_/X _11417_/B VGND VGND VPWR VPWR _11251_/X sky130_fd_sc_hd__o21a_1
X_11182_ _09140_/Y _11181_/A _09140_/A _11181_/Y _09204_/X VGND VGND VPWR VPWR _13367_/A
+ sky130_fd_sc_hd__a221o_2
X_10202_ _09403_/X _08931_/Y _09404_/Y _08931_/A VGND VGND VPWR VPWR _11243_/A sky130_fd_sc_hd__a22o_2
XFILLER_69_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10133_ _10133_/A _10133_/B VGND VGND VPWR VPWR _10134_/B sky130_fd_sc_hd__or2_1
XFILLER_121_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15990_ _15991_/A _15991_/B VGND VGND VPWR VPWR _15992_/A sky130_fd_sc_hd__and2_1
XFILLER_95_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14941_ _14939_/Y _14940_/X _14939_/Y _14940_/X VGND VGND VPWR VPWR _14980_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10064_ _10063_/A _10063_/B _09963_/A _10063_/X VGND VGND VPWR VPWR _10067_/A sky130_fd_sc_hd__a22o_1
X_14872_ _14872_/A VGND VGND VPWR VPWR _15546_/A sky130_fd_sc_hd__buf_1
XFILLER_48_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13823_ _13760_/X _13822_/X _13760_/X _13822_/X VGND VGND VPWR VPWR _13844_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13754_ _13754_/A _13754_/B VGND VGND VPWR VPWR _13755_/A sky130_fd_sc_hd__or2_1
XFILLER_71_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10966_ _10966_/A VGND VGND VPWR VPWR _11604_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16473_ _16473_/D _16454_/Y VGND VGND VPWR VPWR _16473_/Q sky130_fd_sc_hd__dlxtn_1
X_10897_ _10767_/X _10896_/X _10767_/X _10896_/X VGND VGND VPWR VPWR _10909_/B sky130_fd_sc_hd__a2bb2o_1
X_13685_ _13684_/A _13684_/B _11959_/X _13684_/X VGND VGND VPWR VPWR _13686_/A sky130_fd_sc_hd__o22a_1
XFILLER_71_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12705_ _12704_/Y _12656_/Y _12704_/Y _12656_/Y VGND VGND VPWR VPWR _12706_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12636_ _14178_/A _12634_/X _12635_/X VGND VGND VPWR VPWR _12636_/X sky130_fd_sc_hd__o21a_1
X_15424_ _15286_/X _15423_/X _15286_/X _15423_/X VGND VGND VPWR VPWR _15424_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15355_ _15290_/X _15354_/X _15290_/X _15354_/X VGND VGND VPWR VPWR _15422_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14306_ _15966_/A _14396_/B VGND VGND VPWR VPWR _15583_/A sky130_fd_sc_hd__and2_1
X_12567_ _12567_/A VGND VGND VPWR VPWR _12567_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12498_ _12648_/A VGND VGND VPWR VPWR _12499_/A sky130_fd_sc_hd__inv_2
X_15286_ _15287_/A _15284_/Y _15287_/B VGND VGND VPWR VPWR _15286_/X sky130_fd_sc_hd__o21ba_1
X_11518_ _11518_/A _11518_/B VGND VGND VPWR VPWR _11518_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14237_ _14237_/A VGND VGND VPWR VPWR _14243_/A sky130_fd_sc_hd__inv_2
X_11449_ _11449_/A VGND VGND VPWR VPWR _14109_/A sky130_fd_sc_hd__buf_1
XFILLER_50_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14168_ _13448_/A _14145_/A _14143_/Y VGND VGND VPWR VPWR _14168_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13119_ _15243_/A _13119_/B VGND VGND VPWR VPWR _13119_/Y sky130_fd_sc_hd__nand2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _15461_/A _14032_/B _14032_/A _14032_/B VGND VGND VPWR VPWR _14099_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08660_ _08660_/A _08662_/B VGND VGND VPWR VPWR _08919_/A sky130_fd_sc_hd__or2b_1
XFILLER_66_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08591_ _08794_/A _09213_/B _08794_/A _09213_/B VGND VGND VPWR VPWR _08592_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_81_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09212_ _09212_/A VGND VGND VPWR VPWR _09212_/Y sky130_fd_sc_hd__inv_2
X_09143_ _09432_/A _09175_/B VGND VGND VPWR VPWR _09143_/Y sky130_fd_sc_hd__nand2_1
X_09074_ _10015_/B _09074_/B VGND VGND VPWR VPWR _09075_/B sky130_fd_sc_hd__or2_1
XFILLER_131_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09976_ _09971_/Y _09974_/Y _09975_/Y VGND VGND VPWR VPWR _09978_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08927_ _10102_/A _09680_/A VGND VGND VPWR VPWR _08928_/A sky130_fd_sc_hd__or2_2
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08858_ _09502_/A _08842_/Y _08844_/Y _08857_/X VGND VGND VPWR VPWR _08955_/A sky130_fd_sc_hd__o22a_1
XFILLER_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08789_ _08789_/A VGND VGND VPWR VPWR _08789_/Y sky130_fd_sc_hd__inv_2
X_10820_ _10819_/A _10818_/Y _10819_/Y _10818_/A _10974_/A VGND VGND VPWR VPWR _10964_/B
+ sky130_fd_sc_hd__a221o_1
X_10751_ _13757_/A VGND VGND VPWR VPWR _11964_/A sky130_fd_sc_hd__inv_2
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13470_ _13466_/X _13469_/X _13466_/X _13469_/X VGND VGND VPWR VPWR _13470_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12421_ _12432_/B VGND VGND VPWR VPWR _12421_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10682_ _10681_/A _10680_/Y _10681_/Y _10680_/A _10974_/A VGND VGND VPWR VPWR _10811_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12352_ _12309_/A _12309_/B _12309_/Y _12533_/A VGND VGND VPWR VPWR _12525_/A sky130_fd_sc_hd__a2bb2o_1
X_15140_ _15140_/A _15140_/B VGND VGND VPWR VPWR _15140_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12283_ _12258_/X _12282_/Y _12258_/X _12282_/Y VGND VGND VPWR VPWR _12362_/B sky130_fd_sc_hd__a2bb2o_1
X_15071_ _15035_/X _15070_/X _15035_/X _15070_/X VGND VGND VPWR VPWR _15072_/B sky130_fd_sc_hd__a2bb2o_1
X_11303_ _11302_/A _11302_/B _11302_/X _11129_/X VGND VGND VPWR VPWR _11303_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14022_ _15408_/A _13950_/B _13950_/Y VGND VGND VPWR VPWR _14022_/Y sky130_fd_sc_hd__o21ai_1
X_11234_ _11234_/A _11079_/X VGND VGND VPWR VPWR _11234_/X sky130_fd_sc_hd__or2b_1
XFILLER_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11165_ _13716_/A _11295_/B _11164_/Y VGND VGND VPWR VPWR _11165_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15973_ _15993_/A _15971_/X _15972_/X VGND VGND VPWR VPWR _15973_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10116_ _10116_/A _10116_/B VGND VGND VPWR VPWR _10117_/A sky130_fd_sc_hd__or2_1
X_11096_ _11096_/A _11096_/B VGND VGND VPWR VPWR _11096_/Y sky130_fd_sc_hd__nand2_1
X_14924_ _15548_/A _14924_/B VGND VGND VPWR VPWR _14924_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10047_ _10047_/A _10047_/B VGND VGND VPWR VPWR _10047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14855_ _15353_/A _14958_/B _14854_/Y VGND VGND VPWR VPWR _14855_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08231__2 _16357_/A VGND VGND VPWR VPWR _08232_/A sky130_fd_sc_hd__inv_2
X_14786_ _14786_/A _14786_/B VGND VGND VPWR VPWR _14786_/X sky130_fd_sc_hd__and2_1
X_13806_ _14410_/A _13856_/B VGND VGND VPWR VPWR _13806_/Y sky130_fd_sc_hd__nor2_1
X_11998_ _11998_/A _11997_/X VGND VGND VPWR VPWR _11998_/X sky130_fd_sc_hd__or2b_1
XFILLER_16_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13737_ _13694_/X _13736_/X _13694_/X _13736_/X VGND VGND VPWR VPWR _13765_/B sky130_fd_sc_hd__a2bb2o_1
X_10949_ _12940_/A VGND VGND VPWR VPWR _12095_/A sky130_fd_sc_hd__inv_2
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16456_ VGND VGND VPWR VPWR _16456_/HI _16456_/LO sky130_fd_sc_hd__conb_1
X_15407_ _15456_/A _15405_/X _15406_/X VGND VGND VPWR VPWR _15407_/X sky130_fd_sc_hd__o21a_1
X_13668_ _15134_/A _13626_/B _13626_/Y VGND VGND VPWR VPWR _13668_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16387_ _16124_/X _16386_/X _16124_/X _16386_/X VGND VGND VPWR VPWR _16388_/B sky130_fd_sc_hd__a2bb2o_1
X_12619_ _12619_/A _12619_/B VGND VGND VPWR VPWR _12619_/X sky130_fd_sc_hd__or2_1
X_13599_ _13625_/A _13626_/B VGND VGND VPWR VPWR _13599_/Y sky130_fd_sc_hd__nor2_1
X_15338_ _15381_/A _15336_/X _15337_/X VGND VGND VPWR VPWR _15338_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_0 _12648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15269_ _15212_/X _15268_/X _15212_/X _15268_/X VGND VGND VPWR VPWR _15270_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _09830_/A VGND VGND VPWR VPWR _09830_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09736_/A _09736_/B _09739_/A VGND VGND VPWR VPWR _10046_/A sky130_fd_sc_hd__a21bo_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08712_/A _09470_/B VGND VGND VPWR VPWR _08712_/Y sky130_fd_sc_hd__nor2_1
X_09692_ _09692_/A _09692_/B VGND VGND VPWR VPWR _09695_/A sky130_fd_sc_hd__or2_1
Xrebuffer12 rebuffer13/X VGND VGND VPWR VPWR rebuffer12/X sky130_fd_sc_hd__dlygate4sd1_1
X_08643_ _08718_/A VGND VGND VPWR VPWR _09458_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer34 _08358_/A VGND VGND VPWR VPWR _08281_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer23 _10194_/B VGND VGND VPWR VPWR rebuffer23/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08574_ _08574_/A VGND VGND VPWR VPWR _08574_/Y sky130_fd_sc_hd__inv_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09126_ _09701_/A _09126_/B VGND VGND VPWR VPWR _09126_/Y sky130_fd_sc_hd__nand2_1
X_09057_ _08789_/Y _09050_/A _08789_/A _09050_/Y VGND VGND VPWR VPWR _10013_/B sky130_fd_sc_hd__o22a_1
XFILLER_116_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09959_ _09951_/Y _09957_/Y _09958_/Y VGND VGND VPWR VPWR _09972_/B sky130_fd_sc_hd__o21ai_1
XFILLER_131_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12970_ _13701_/A VGND VGND VPWR VPWR _14524_/A sky130_fd_sc_hd__inv_2
XFILLER_18_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11921_ _10559_/A _11856_/A _10673_/B _11920_/Y VGND VGND VPWR VPWR _11922_/A sky130_fd_sc_hd__o22a_1
X_14640_ _14573_/X _14639_/Y _14573_/X _14639_/Y VGND VGND VPWR VPWR _14646_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11852_ _11852_/A _11852_/B VGND VGND VPWR VPWR _11852_/X sky130_fd_sc_hd__or2_1
X_14571_ _15270_/A _14572_/B VGND VGND VPWR VPWR _14571_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10803_ _09987_/A _09987_/B _09987_/Y VGND VGND VPWR VPWR _10804_/A sky130_fd_sc_hd__o21ai_1
X_16310_ _16250_/X _16309_/Y _16250_/X _16309_/Y VGND VGND VPWR VPWR _16318_/B sky130_fd_sc_hd__o2bb2a_1
X_11783_ _11783_/A _11784_/B VGND VGND VPWR VPWR _11785_/A sky130_fd_sc_hd__and2_1
X_13522_ _13522_/A _13522_/B VGND VGND VPWR VPWR _13522_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10734_ _11968_/A VGND VGND VPWR VPWR _13083_/A sky130_fd_sc_hd__buf_1
X_16241_ _16241_/A VGND VGND VPWR VPWR _16241_/Y sky130_fd_sc_hd__inv_2
X_13453_ _13452_/Y _13307_/X _13209_/Y VGND VGND VPWR VPWR _13453_/Y sky130_fd_sc_hd__o21ai_1
X_10665_ _09984_/A _09984_/B _09984_/Y VGND VGND VPWR VPWR _10666_/A sky130_fd_sc_hd__o21ai_1
X_16172_ _16109_/X _16171_/X _16109_/X _16171_/X VGND VGND VPWR VPWR _16173_/B sky130_fd_sc_hd__a2bb2oi_1
X_13384_ _14132_/A _13444_/B VGND VGND VPWR VPWR _13384_/Y sky130_fd_sc_hd__nor2_1
X_12404_ _12404_/A _12404_/B VGND VGND VPWR VPWR _12404_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12335_ _12331_/Y _12580_/A _12334_/Y VGND VGND VPWR VPWR _12339_/B sky130_fd_sc_hd__o21ai_1
X_15123_ _15066_/A _15066_/B _15066_/Y VGND VGND VPWR VPWR _15123_/Y sky130_fd_sc_hd__o21ai_1
X_10596_ _10596_/A VGND VGND VPWR VPWR _10596_/Y sky130_fd_sc_hd__inv_2
X_15054_ _15054_/A _15054_/B VGND VGND VPWR VPWR _15054_/Y sky130_fd_sc_hd__nand2_1
X_12266_ _12266_/A _12266_/B VGND VGND VPWR VPWR _12266_/X sky130_fd_sc_hd__or2_1
XFILLER_5_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14005_ _13961_/X _14004_/Y _13961_/X _14004_/Y VGND VGND VPWR VPWR _14066_/B sky130_fd_sc_hd__a2bb2o_1
X_11217_ _11084_/X _11216_/X _11084_/X _11216_/X VGND VGND VPWR VPWR _11218_/B sky130_fd_sc_hd__a2bb2o_1
X_12197_ _13202_/A _12249_/B _12196_/Y VGND VGND VPWR VPWR _12197_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11148_ _11148_/A VGND VGND VPWR VPWR _11148_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15956_ _15956_/A _15956_/B VGND VGND VPWR VPWR _15956_/X sky130_fd_sc_hd__or2_1
X_11079_ _13926_/A _11079_/B VGND VGND VPWR VPWR _11079_/X sky130_fd_sc_hd__or2_1
XFILLER_49_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15887_ _15883_/Y _15885_/X _15886_/Y VGND VGND VPWR VPWR _15887_/X sky130_fd_sc_hd__o21a_1
X_14907_ _14901_/Y _14905_/X _14906_/Y VGND VGND VPWR VPWR _14907_/X sky130_fd_sc_hd__o21a_1
X_14838_ _14754_/A _14754_/B _14751_/X _14754_/Y VGND VGND VPWR VPWR _14838_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14769_ _14744_/X _14768_/Y _14744_/X _14768_/Y VGND VGND VPWR VPWR _14771_/B sky130_fd_sc_hd__a2bb2o_1
X_08290_ _08331_/A input32/X _08332_/A _08334_/A VGND VGND VPWR VPWR _08329_/A sky130_fd_sc_hd__o22a_1
XFILLER_32_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16439_ _16419_/B _16436_/X _16435_/X _16438_/X VGND VGND VPWR VPWR _16439_/X sky130_fd_sc_hd__o22a_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09813_ _09812_/X _08813_/A _09812_/X _08813_/A VGND VGND VPWR VPWR _09821_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09744_ _08524_/Y _09743_/X _08524_/Y _09743_/X VGND VGND VPWR VPWR _09745_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09675_ _10930_/A _09675_/B VGND VGND VPWR VPWR _11939_/A sky130_fd_sc_hd__or2_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08626_ _08625_/A _08365_/Y _08625_/Y _08365_/A VGND VGND VPWR VPWR _08627_/B sky130_fd_sc_hd__o22a_1
XFILLER_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08557_ _09737_/A _08567_/B VGND VGND VPWR VPWR _08558_/A sky130_fd_sc_hd__or2_1
X_08488_ _08263_/A _08341_/B _08476_/Y _08587_/A VGND VGND VPWR VPWR _08574_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10450_ _11803_/A VGND VGND VPWR VPWR _11764_/A sky130_fd_sc_hd__inv_2
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09109_ _09714_/A _09107_/B _09107_/X _09108_/Y VGND VGND VPWR VPWR _09113_/B sky130_fd_sc_hd__o22ai_2
X_10381_ _10381_/A VGND VGND VPWR VPWR _10381_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12120_ _13190_/A _12055_/B _12055_/Y VGND VGND VPWR VPWR _12120_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12051_ _12051_/A _12051_/B VGND VGND VPWR VPWR _12051_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11002_ _11002_/A VGND VGND VPWR VPWR _14410_/A sky130_fd_sc_hd__buf_1
XFILLER_77_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15810_ _15749_/Y _15808_/X _15809_/Y VGND VGND VPWR VPWR _15810_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15741_ _15679_/A _15679_/B _15679_/Y VGND VGND VPWR VPWR _15741_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12953_ _12953_/A VGND VGND VPWR VPWR _13879_/A sky130_fd_sc_hd__inv_2
XFILLER_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15672_ _15638_/Y _15670_/X _15671_/Y VGND VGND VPWR VPWR _15672_/X sky130_fd_sc_hd__o21a_1
X_11904_ _11904_/A _11904_/B VGND VGND VPWR VPWR _11904_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14623_ _14623_/A VGND VGND VPWR VPWR _15339_/A sky130_fd_sc_hd__buf_1
X_12884_ _12936_/A VGND VGND VPWR VPWR _14477_/A sky130_fd_sc_hd__buf_1
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11835_/A _11835_/B VGND VGND VPWR VPWR _11835_/Y sky130_fd_sc_hd__nand2_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14515_/X _14553_/X _14515_/X _14553_/X VGND VGND VPWR VPWR _14580_/B sky130_fd_sc_hd__a2bb2o_1
X_11766_ _11803_/B _11765_/X _11803_/B _11765_/X VGND VGND VPWR VPWR _11799_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _14485_/A VGND VGND VPWR VPWR _15199_/A sky130_fd_sc_hd__buf_1
X_10717_ _11904_/A VGND VGND VPWR VPWR _13695_/A sky130_fd_sc_hd__buf_1
X_13505_ _13507_/A VGND VGND VPWR VPWR _15044_/A sky130_fd_sc_hd__buf_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16224_ _16224_/A VGND VGND VPWR VPWR _16224_/Y sky130_fd_sc_hd__inv_2
X_13436_ _14112_/A _13436_/B VGND VGND VPWR VPWR _13436_/Y sky130_fd_sc_hd__nand2_1
X_11697_ _11637_/A _11639_/X _11636_/X VGND VGND VPWR VPWR _11697_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer3 _08361_/A VGND VGND VPWR VPWR _08404_/B1 sky130_fd_sc_hd__dlygate4sd1_1
X_10648_ _09969_/Y _10647_/A _10077_/A _10647_/Y _10940_/A VGND VGND VPWR VPWR _11978_/A
+ sky130_fd_sc_hd__a221o_2
X_16155_ _16067_/X _16155_/B VGND VGND VPWR VPWR _16155_/X sky130_fd_sc_hd__and2b_1
X_13367_ _13367_/A _13367_/B VGND VGND VPWR VPWR _13367_/X sky130_fd_sc_hd__or2_1
X_10579_ _11867_/A _10651_/B VGND VGND VPWR VPWR _10579_/Y sky130_fd_sc_hd__nand2_1
X_16086_ _16089_/A _16089_/B VGND VGND VPWR VPWR _16086_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12318_ _14082_/A _12318_/B VGND VGND VPWR VPWR _12319_/A sky130_fd_sc_hd__nand2_1
X_13298_ _13230_/Y _13296_/Y _13297_/Y VGND VGND VPWR VPWR _13299_/A sky130_fd_sc_hd__o21ai_2
X_15106_ _15100_/X _15105_/X _15100_/X _15105_/X VGND VGND VPWR VPWR _15107_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12249_ _13202_/A _12249_/B VGND VGND VPWR VPWR _12249_/Y sky130_fd_sc_hd__nor2_1
X_15037_ _15070_/A _15035_/X _15036_/X VGND VGND VPWR VPWR _15037_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15939_ _15952_/A _15952_/B VGND VGND VPWR VPWR _16017_/A sky130_fd_sc_hd__and2_1
XFILLER_37_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09460_ _09460_/A VGND VGND VPWR VPWR _09460_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08411_ _09225_/A VGND VGND VPWR VPWR _08717_/A sky130_fd_sc_hd__inv_2
X_09391_ _10420_/B VGND VGND VPWR VPWR _09392_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08342_ _08342_/A _08342_/B VGND VGND VPWR VPWR _08343_/A sky130_fd_sc_hd__or2_1
X_08273_ input10/X VGND VGND VPWR VPWR _08357_/B sky130_fd_sc_hd__inv_2
XFILLER_20_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09727_ _09727_/A VGND VGND VPWR VPWR _09727_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09658_ _09987_/A _09658_/B VGND VGND VPWR VPWR _09658_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _08229_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_82_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08609_ _08609_/A VGND VGND VPWR VPWR _10113_/B sky130_fd_sc_hd__inv_2
X_09589_ _08688_/A _09019_/A _09532_/A VGND VGND VPWR VPWR _09589_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11620_/A _12379_/A VGND VGND VPWR VPWR _11620_/Y sky130_fd_sc_hd__nor2_1
X_11551_ _11486_/Y _11550_/Y _11486_/Y _11550_/Y VGND VGND VPWR VPWR _11554_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10502_ _12926_/A VGND VGND VPWR VPWR _11837_/A sky130_fd_sc_hd__inv_2
X_14270_ _14198_/Y _14268_/Y _14269_/Y VGND VGND VPWR VPWR _14271_/A sky130_fd_sc_hd__o21ai_2
XFILLER_109_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11482_ _09788_/A _09368_/A _09430_/X VGND VGND VPWR VPWR _11482_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13221_ _15057_/A VGND VGND VPWR VPWR _14674_/A sky130_fd_sc_hd__inv_2
X_10433_ _10512_/A _10431_/X _10432_/X VGND VGND VPWR VPWR _10433_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13152_ _13118_/X _13151_/Y _13118_/X _13151_/Y VGND VGND VPWR VPWR _13200_/B sky130_fd_sc_hd__a2bb2o_1
X_10364_ _11755_/A VGND VGND VPWR VPWR _13522_/A sky130_fd_sc_hd__buf_1
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12103_ _12067_/X _12102_/Y _12067_/X _12102_/Y VGND VGND VPWR VPWR _12155_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13083_ _13083_/A VGND VGND VPWR VPWR _13761_/A sky130_fd_sc_hd__inv_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _12706_/A _10291_/B _10291_/X _10294_/Y VGND VGND VPWR VPWR _10295_/X sky130_fd_sc_hd__a22o_1
X_12034_ _13188_/A _12053_/B VGND VGND VPWR VPWR _12034_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13985_ _13985_/A _13985_/B VGND VGND VPWR VPWR _13985_/X sky130_fd_sc_hd__or2_1
XFILLER_46_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15724_ _15684_/X _15723_/Y _15684_/X _15723_/Y VGND VGND VPWR VPWR _15817_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12936_ _12936_/A _12936_/B VGND VGND VPWR VPWR _12936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15655_ _15778_/A _15655_/B VGND VGND VPWR VPWR _15656_/A sky130_fd_sc_hd__or2_1
XFILLER_61_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12867_ _12946_/A _12947_/B VGND VGND VPWR VPWR _12867_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15586_ _15500_/X _15586_/B VGND VGND VPWR VPWR _15586_/X sky130_fd_sc_hd__and2b_1
X_14606_ _14591_/X _14605_/X _14591_/X _14605_/X VGND VGND VPWR VPWR _14665_/B sky130_fd_sc_hd__a2bb2o_1
X_11818_ _13629_/A _11843_/B VGND VGND VPWR VPWR _11818_/Y sky130_fd_sc_hd__nor2_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14537_/A _14536_/X VGND VGND VPWR VPWR _14537_/X sky130_fd_sc_hd__or2b_1
X_12798_ _12856_/A _12856_/B VGND VGND VPWR VPWR _12798_/Y sky130_fd_sc_hd__nor2_1
X_11749_ _11750_/A _11750_/B VGND VGND VPWR VPWR _11751_/A sky130_fd_sc_hd__and2_1
X_14468_ _14445_/Y _14466_/X _14467_/Y VGND VGND VPWR VPWR _14468_/X sky130_fd_sc_hd__o21a_1
X_16207_ _16207_/A VGND VGND VPWR VPWR _16207_/Y sky130_fd_sc_hd__inv_2
X_14399_ _14399_/A _14286_/X VGND VGND VPWR VPWR _14399_/X sky130_fd_sc_hd__or2b_1
X_13419_ _13340_/A _13340_/B _13340_/A _13340_/B VGND VGND VPWR VPWR _13419_/X sky130_fd_sc_hd__a2bb2o_1
X_16138_ _16138_/A _16121_/X VGND VGND VPWR VPWR _16139_/A sky130_fd_sc_hd__or2b_1
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16069_ _16043_/X _16068_/Y _16043_/X _16068_/Y VGND VGND VPWR VPWR _16112_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08960_ _08960_/A _08960_/B VGND VGND VPWR VPWR _08960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08891_ _09555_/A _08571_/A _08573_/A VGND VGND VPWR VPWR _08891_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09512_ _08795_/X _09492_/B _09492_/Y _09511_/X VGND VGND VPWR VPWR _09512_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09443_ _09441_/X _09442_/X _09441_/X _09442_/X VGND VGND VPWR VPWR _10904_/A sky130_fd_sc_hd__a2bb2oi_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09374_ _09374_/A VGND VGND VPWR VPWR _09431_/B sky130_fd_sc_hd__inv_2
X_08325_ _08323_/Y _08324_/A _08323_/A _08324_/Y _08304_/X VGND VGND VPWR VPWR _08555_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08256_ input32/X VGND VGND VPWR VPWR _08257_/B sky130_fd_sc_hd__inv_2
XFILLER_106_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10080_ _10049_/X _10078_/X _10813_/B VGND VGND VPWR VPWR _10080_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13770_ _13810_/A _13768_/X _13769_/X VGND VGND VPWR VPWR _13770_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10982_ _10982_/A VGND VGND VPWR VPWR _10982_/X sky130_fd_sc_hd__clkbuf_2
X_12721_ _12680_/X _12720_/X _12680_/X _12720_/X VGND VGND VPWR VPWR _13458_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15440_ _15440_/A _15440_/B VGND VGND VPWR VPWR _15440_/X sky130_fd_sc_hd__and2_1
X_12652_ _15285_/A VGND VGND VPWR VPWR _13985_/A sky130_fd_sc_hd__inv_2
XFILLER_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11603_ _10088_/X _11602_/X _10088_/X _11602_/X VGND VGND VPWR VPWR _11604_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12583_ _12580_/Y _12582_/Y _12580_/A _12582_/A _12500_/A VGND VGND VPWR VPWR _12621_/B
+ sky130_fd_sc_hd__o221a_1
X_15371_ _15412_/A _15412_/B VGND VGND VPWR VPWR _15447_/A sky130_fd_sc_hd__and2_1
XFILLER_129_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14322_ _15863_/A _14269_/B _14269_/Y VGND VGND VPWR VPWR _14322_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11534_ _11533_/A _11533_/B _11533_/Y _10982_/X VGND VGND VPWR VPWR _12416_/A sky130_fd_sc_hd__o211a_2
XFILLER_128_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14253_ _14253_/A VGND VGND VPWR VPWR _14253_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11465_ _14064_/A VGND VGND VPWR VPWR _15440_/A sky130_fd_sc_hd__buf_1
XFILLER_7_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13204_ _13204_/A _13204_/B VGND VGND VPWR VPWR _13204_/Y sky130_fd_sc_hd__nand2_1
X_10416_ _08402_/X _10277_/A _08929_/A _10339_/Y _10420_/B VGND VGND VPWR VPWR _10429_/A
+ sky130_fd_sc_hd__o221a_1
X_14184_ _14184_/A _12633_/X VGND VGND VPWR VPWR _14184_/X sky130_fd_sc_hd__or2b_1
X_11396_ _11393_/Y _11395_/Y _11393_/A _11395_/A _12605_/B VGND VGND VPWR VPWR _13396_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_124_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13135_ _15167_/A VGND VGND VPWR VPWR _14934_/A sky130_fd_sc_hd__clkbuf_2
X_10347_ _10347_/A VGND VGND VPWR VPWR _11711_/B sky130_fd_sc_hd__inv_2
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _13023_/X _13065_/X _13023_/X _13065_/X VGND VGND VPWR VPWR _13115_/B sky130_fd_sc_hd__a2bb2o_1
X_10278_ _08929_/A _10277_/A _08402_/X _10277_/Y _10268_/A VGND VGND VPWR VPWR _11713_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_3_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12017_ _11975_/X _12016_/Y _11975_/X _12016_/Y VGND VGND VPWR VPWR _12061_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13968_ _15167_/A _13968_/B VGND VGND VPWR VPWR _13968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15707_ _15552_/A _14928_/B _14928_/Y VGND VGND VPWR VPWR _15707_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12919_ _12919_/A VGND VGND VPWR VPWR _13002_/A sky130_fd_sc_hd__inv_2
XFILLER_46_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13899_ _14410_/A _13856_/B _13856_/Y VGND VGND VPWR VPWR _13899_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15638_ _15671_/A _15671_/B VGND VGND VPWR VPWR _15638_/Y sky130_fd_sc_hd__nor2_1
X_15569_ _15429_/X _15568_/X _15429_/X _15568_/X VGND VGND VPWR VPWR _15655_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09090_ _09701_/A VGND VGND VPWR VPWR _09421_/A sky130_fd_sc_hd__buf_1
XFILLER_115_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09992_ _09992_/A _09993_/B VGND VGND VPWR VPWR _09992_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08943_ _08939_/Y _11405_/A _08942_/Y VGND VGND VPWR VPWR _08952_/A sky130_fd_sc_hd__o21ai_2
XFILLER_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08874_ _08873_/Y _08867_/X _08873_/Y _08867_/X VGND VGND VPWR VPWR _08984_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09426_ _09426_/A _09433_/B VGND VGND VPWR VPWR _09426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09357_ _08692_/A _09861_/A _09351_/Y _09356_/X VGND VGND VPWR VPWR _09357_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08308_ _08308_/A VGND VGND VPWR VPWR _08308_/Y sky130_fd_sc_hd__inv_2
X_09288_ _09230_/A _09800_/A _09230_/Y VGND VGND VPWR VPWR _09288_/Y sky130_fd_sc_hd__a21oi_1
X_08239_ _08239_/A VGND VGND VPWR VPWR _08239_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11250_ _14048_/A _11250_/B VGND VGND VPWR VPWR _11417_/B sky130_fd_sc_hd__or2_1
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10201_ _10213_/A _10213_/B VGND VGND VPWR VPWR _10201_/Y sky130_fd_sc_hd__nor2_1
X_11181_ _11181_/A VGND VGND VPWR VPWR _11181_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10132_ _10132_/A _10132_/B VGND VGND VPWR VPWR _10133_/B sky130_fd_sc_hd__or2_1
XFILLER_121_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14940_ _14841_/A _14841_/B _14838_/X _14841_/Y VGND VGND VPWR VPWR _14940_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10063_ _10063_/A _10063_/B VGND VGND VPWR VPWR _10063_/X sky130_fd_sc_hd__or2_1
X_14871_ _15548_/A _14924_/B VGND VGND VPWR VPWR _14871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13822_ _13822_/A _13761_/X VGND VGND VPWR VPWR _13822_/X sky130_fd_sc_hd__or2b_1
XFILLER_75_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13753_ _13753_/A _13753_/B VGND VGND VPWR VPWR _13753_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12704_ _12704_/A VGND VGND VPWR VPWR _12704_/Y sky130_fd_sc_hd__inv_2
X_10965_ _10964_/Y _10812_/X _10821_/Y VGND VGND VPWR VPWR _10965_/X sky130_fd_sc_hd__o21a_1
X_16472_ _16472_/D _16456_/LO VGND VGND VPWR VPWR _16472_/Q sky130_fd_sc_hd__dlxtn_1
X_10896_ _10896_/A _10769_/X VGND VGND VPWR VPWR _10896_/X sky130_fd_sc_hd__or2b_1
X_13684_ _13684_/A _13684_/B VGND VGND VPWR VPWR _13684_/X sky130_fd_sc_hd__and2_1
X_12635_ _12635_/A _12635_/B VGND VGND VPWR VPWR _12635_/X sky130_fd_sc_hd__or2_1
XFILLER_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15423_ _15356_/Y _15421_/Y _15422_/Y VGND VGND VPWR VPWR _15423_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12566_ _14912_/A _11440_/B _11440_/Y VGND VGND VPWR VPWR _12567_/A sky130_fd_sc_hd__o21ai_1
X_15354_ _15357_/A _15352_/X _15353_/X VGND VGND VPWR VPWR _15354_/X sky130_fd_sc_hd__o21a_1
X_14305_ _14277_/A _14304_/Y _14277_/A _14304_/Y VGND VGND VPWR VPWR _14396_/B sky130_fd_sc_hd__a2bb2o_1
X_11517_ _11513_/Y _12684_/A _11313_/X _11516_/Y VGND VGND VPWR VPWR _11517_/X sky130_fd_sc_hd__o22a_1
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12497_ _12473_/X _12496_/X _12473_/X _12496_/X VGND VGND VPWR VPWR _12648_/A sky130_fd_sc_hd__a2bb2o_4
X_15285_ _15285_/A _15285_/B VGND VGND VPWR VPWR _15287_/B sky130_fd_sc_hd__and2_1
X_14236_ _14236_/A _15839_/A VGND VGND VPWR VPWR _14237_/A sky130_fd_sc_hd__or2_1
X_11448_ _12349_/A _11453_/B VGND VGND VPWR VPWR _11448_/Y sky130_fd_sc_hd__nor2_1
X_14167_ _14167_/A _14166_/X VGND VGND VPWR VPWR _14167_/X sky130_fd_sc_hd__or2b_1
X_11379_ _08973_/X _11378_/X _08973_/X _11378_/X VGND VGND VPWR VPWR _11380_/B sky130_fd_sc_hd__a2bb2oi_2
X_13118_ _13062_/Y _13116_/X _13117_/Y VGND VGND VPWR VPWR _13118_/X sky130_fd_sc_hd__o21a_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14098_/A _14101_/B VGND VGND VPWR VPWR _14098_/Y sky130_fd_sc_hd__nor2_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13049_ _13775_/A VGND VGND VPWR VPWR _15240_/A sky130_fd_sc_hd__buf_1
XFILLER_66_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08590_ _09455_/B VGND VGND VPWR VPWR _09551_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09211_ _09553_/A _09731_/A VGND VGND VPWR VPWR _09212_/A sky130_fd_sc_hd__or2_1
X_09142_ _09138_/Y _09140_/Y _09141_/Y VGND VGND VPWR VPWR _09175_/B sky130_fd_sc_hd__o21ai_1
X_09073_ _10016_/B _09073_/B VGND VGND VPWR VPWR _09074_/B sky130_fd_sc_hd__or2_1
XFILLER_107_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09975_ _09975_/A _09975_/B VGND VGND VPWR VPWR _09975_/Y sky130_fd_sc_hd__nand2_1
X_08926_ _09817_/A VGND VGND VPWR VPWR _10102_/A sky130_fd_sc_hd__inv_2
XFILLER_85_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08857_ _10103_/A _08855_/Y _08916_/A _09460_/A VGND VGND VPWR VPWR _08857_/X sky130_fd_sc_hd__o22a_1
XFILLER_17_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08788_ _08712_/A _09470_/B _08712_/Y VGND VGND VPWR VPWR _08789_/A sky130_fd_sc_hd__a21oi_2
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10750_ _09635_/A _10749_/A _09635_/Y _10749_/Y _09672_/A VGND VGND VPWR VPWR _13757_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_111_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10681_ _10681_/A VGND VGND VPWR VPWR _10681_/Y sky130_fd_sc_hd__inv_2
X_09409_ _09409_/A _09409_/B VGND VGND VPWR VPWR _09409_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12420_ _12419_/A _12419_/B _12419_/Y VGND VGND VPWR VPWR _12432_/B sky130_fd_sc_hd__o21ai_2
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12351_ _12312_/A _12312_/B _12312_/Y _12541_/A VGND VGND VPWR VPWR _12533_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12282_ _13789_/A _12365_/B _12281_/Y VGND VGND VPWR VPWR _12282_/Y sky130_fd_sc_hd__o21ai_1
X_15070_ _15070_/A _15036_/X VGND VGND VPWR VPWR _15070_/X sky130_fd_sc_hd__or2b_1
X_11302_ _11302_/A _11302_/B VGND VGND VPWR VPWR _11302_/X sky130_fd_sc_hd__and2_1
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11233_ _12227_/A VGND VGND VPWR VPWR _13341_/A sky130_fd_sc_hd__buf_1
X_14021_ _14021_/A _14056_/B VGND VGND VPWR VPWR _14077_/A sky130_fd_sc_hd__and2_1
XFILLER_5_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11164_ _12187_/A _11295_/B VGND VGND VPWR VPWR _11164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15972_ _15972_/A _15972_/B VGND VGND VPWR VPWR _15972_/X sky130_fd_sc_hd__or2_1
XFILLER_95_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10115_ _10115_/A _10115_/B VGND VGND VPWR VPWR _10116_/A sky130_fd_sc_hd__or2_1
X_11095_ _09432_/B _09383_/B _09383_/X VGND VGND VPWR VPWR _11096_/B sky130_fd_sc_hd__a21boi_1
X_14923_ _14875_/Y _14921_/X _14922_/Y VGND VGND VPWR VPWR _14923_/X sky130_fd_sc_hd__o21a_1
X_10046_ _10046_/A _10081_/B VGND VGND VPWR VPWR _10046_/X sky130_fd_sc_hd__and2_1
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14854_ _15353_/A _14958_/B VGND VGND VPWR VPWR _14854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14785_ _14736_/X _14784_/X _14736_/X _14784_/X VGND VGND VPWR VPWR _14786_/B sky130_fd_sc_hd__a2bb2o_1
X_13805_ _13772_/X _13804_/X _13772_/X _13804_/X VGND VGND VPWR VPWR _13856_/B sky130_fd_sc_hd__a2bb2o_1
X_11997_ _11997_/A _11997_/B VGND VGND VPWR VPWR _11997_/X sky130_fd_sc_hd__or2_1
X_13736_ _13736_/A _13695_/X VGND VGND VPWR VPWR _13736_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10948_ _10946_/Y _10947_/Y _10947_/B _09916_/X _10792_/X VGND VGND VPWR VPWR _12940_/A
+ sky130_fd_sc_hd__o221a_2
X_16455_ _16471_/Q _08230_/A _08233_/A _16392_/C _16343_/A VGND VGND VPWR VPWR _16471_/D
+ sky130_fd_sc_hd__o221a_2
X_15406_ _15406_/A _15406_/B VGND VGND VPWR VPWR _15406_/X sky130_fd_sc_hd__or2_1
X_10879_ _12053_/A VGND VGND VPWR VPWR _10883_/A sky130_fd_sc_hd__inv_2
X_13667_ _13695_/A _13695_/B VGND VGND VPWR VPWR _13736_/A sky130_fd_sc_hd__and2_1
XFILLER_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16386_ _16058_/X _16386_/B VGND VGND VPWR VPWR _16386_/X sky130_fd_sc_hd__and2b_1
X_12618_ _12604_/X _14236_/A _14232_/B VGND VGND VPWR VPWR _12618_/X sky130_fd_sc_hd__o21a_1
X_13598_ _13577_/X _13597_/Y _13577_/X _13597_/Y VGND VGND VPWR VPWR _13626_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12549_ _12549_/A VGND VGND VPWR VPWR _12549_/Y sky130_fd_sc_hd__inv_2
X_15337_ _15337_/A _15337_/B VGND VGND VPWR VPWR _15337_/X sky130_fd_sc_hd__or2_1
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15268_ _15268_/A _15216_/X VGND VGND VPWR VPWR _15268_/X sky130_fd_sc_hd__or2b_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 input20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14219_ _14231_/A _14219_/B VGND VGND VPWR VPWR _15875_/A sky130_fd_sc_hd__or2_1
XFILLER_125_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15199_ _15199_/A _15199_/B VGND VGND VPWR VPWR _15199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _09760_/A VGND VGND VPWR VPWR _09782_/A sky130_fd_sc_hd__inv_2
XFILLER_79_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _08711_/A _09472_/B VGND VGND VPWR VPWR _08711_/Y sky130_fd_sc_hd__nor2_1
X_09691_ _08618_/X _09693_/B _08618_/X _09693_/B VGND VGND VPWR VPWR _09692_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08642_ _08642_/A VGND VGND VPWR VPWR _08718_/A sky130_fd_sc_hd__inv_2
XFILLER_66_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer24 _10191_/X VGND VGND VPWR VPWR rebuffer24/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer13 rebuffer14/X VGND VGND VPWR VPWR rebuffer13/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08573_ _08573_/A VGND VGND VPWR VPWR _08573_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09125_ _09421_/A _09126_/B VGND VGND VPWR VPWR _09125_/Y sky130_fd_sc_hd__nor2_1
X_09056_ _08781_/Y _09052_/A _08781_/A _09052_/Y VGND VGND VPWR VPWR _10012_/B sky130_fd_sc_hd__o22a_1
XFILLER_89_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09958_ _09958_/A _09958_/B VGND VGND VPWR VPWR _09958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08909_ _08683_/X _08908_/X _08683_/X _08908_/X VGND VGND VPWR VPWR _08970_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09889_ _09874_/X _09888_/X _09874_/X _09888_/X VGND VGND VPWR VPWR _09932_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11920_ _11920_/A _11920_/B VGND VGND VPWR VPWR _11920_/Y sky130_fd_sc_hd__nor2_1
X_11851_ _11913_/A VGND VGND VPWR VPWR _12773_/A sky130_fd_sc_hd__buf_1
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14570_ _13007_/A _14569_/Y _13007_/A _14569_/Y VGND VGND VPWR VPWR _14572_/B sky130_fd_sc_hd__a2bb2o_1
X_11782_ _11787_/A VGND VGND VPWR VPWR _14429_/A sky130_fd_sc_hd__buf_1
X_10802_ _13513_/A _10801_/B _10801_/X _10664_/X VGND VGND VPWR VPWR _10802_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13521_ _10388_/X _13484_/X _10388_/X _13484_/X VGND VGND VPWR VPWR _13522_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10733_ _10731_/A _10732_/A _10731_/Y _10732_/Y _09672_/A VGND VGND VPWR VPWR _11968_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_13_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16240_ _16249_/A _16240_/B VGND VGND VPWR VPWR _16240_/Y sky130_fd_sc_hd__nor2_1
X_13452_ _14934_/A _13452_/B VGND VGND VPWR VPWR _13452_/Y sky130_fd_sc_hd__nor2_1
X_10664_ _13516_/A _10663_/B _10663_/X _10545_/X VGND VGND VPWR VPWR _10664_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16171_ _16073_/X _16171_/B VGND VGND VPWR VPWR _16171_/X sky130_fd_sc_hd__and2b_1
X_13383_ _13368_/X _13382_/X _13368_/X _13382_/X VGND VGND VPWR VPWR _13444_/B sky130_fd_sc_hd__a2bb2o_1
X_12403_ _12357_/X _12402_/X _12357_/X _12402_/X VGND VGND VPWR VPWR _12404_/B sky130_fd_sc_hd__a2bb2o_1
X_10595_ _10595_/A _09717_/X VGND VGND VPWR VPWR _10596_/A sky130_fd_sc_hd__or2b_1
XFILLER_126_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12334_ _12575_/A _12334_/B VGND VGND VPWR VPWR _12334_/Y sky130_fd_sc_hd__nand2_1
X_15122_ _15122_/A _15122_/B VGND VGND VPWR VPWR _15122_/Y sky130_fd_sc_hd__nand2_1
X_15053_ _15047_/X _15052_/X _15047_/X _15052_/X VGND VGND VPWR VPWR _15054_/B sky130_fd_sc_hd__a2bb2o_1
X_14004_ _15420_/A _13962_/B _13962_/Y VGND VGND VPWR VPWR _14004_/Y sky130_fd_sc_hd__o21ai_1
X_12265_ _12369_/A VGND VGND VPWR VPWR _12783_/A sky130_fd_sc_hd__buf_1
X_11216_ _11216_/A _11085_/X VGND VGND VPWR VPWR _11216_/X sky130_fd_sc_hd__or2b_1
X_12196_ _12196_/A _12249_/B VGND VGND VPWR VPWR _12196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11147_ _11147_/A VGND VGND VPWR VPWR _11147_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15955_ _16014_/A _15953_/X _15954_/X VGND VGND VPWR VPWR _15955_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11078_ _14427_/A VGND VGND VPWR VPWR _13926_/A sky130_fd_sc_hd__clkbuf_2
X_15886_ _15886_/A _15886_/B VGND VGND VPWR VPWR _15886_/Y sky130_fd_sc_hd__nand2_1
X_14906_ _14906_/A _14906_/B VGND VGND VPWR VPWR _14906_/Y sky130_fd_sc_hd__nand2_1
X_10029_ _09332_/A _08770_/B _10038_/B _10028_/X VGND VGND VPWR VPWR _10029_/X sky130_fd_sc_hd__o22a_1
X_14837_ _14757_/A _14757_/B _14750_/X _14757_/Y VGND VGND VPWR VPWR _14837_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14768_ _15351_/A _14830_/B _14767_/Y VGND VGND VPWR VPWR _14768_/Y sky130_fd_sc_hd__o21ai_1
X_14699_ _14735_/A _14735_/B VGND VGND VPWR VPWR _14788_/A sky130_fd_sc_hd__and2_1
X_13719_ _13720_/A _13720_/B VGND VGND VPWR VPWR _13721_/A sky130_fd_sc_hd__and2_1
XFILLER_32_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16438_ _16460_/Q _16459_/Q _16458_/Q _16447_/B _16437_/X VGND VGND VPWR VPWR _16438_/X
+ sky130_fd_sc_hd__o41a_1
X_16369_ _16324_/A _16324_/B _16324_/Y VGND VGND VPWR VPWR _16369_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09812_ _08819_/A _08610_/A _09456_/Y _09811_/X VGND VGND VPWR VPWR _09812_/X sky130_fd_sc_hd__o22a_1
XFILLER_101_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09743_ _09743_/A _09743_/B VGND VGND VPWR VPWR _09743_/X sky130_fd_sc_hd__or2_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09674_ _09655_/X _09673_/X _09655_/X _09673_/X VGND VGND VPWR VPWR _09675_/B sky130_fd_sc_hd__a2bb2oi_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08625_ _08625_/A VGND VGND VPWR VPWR _08625_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _16357_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_82_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _09859_/A VGND VGND VPWR VPWR _09737_/A sky130_fd_sc_hd__inv_2
XFILLER_70_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08487_ _08266_/A _08346_/B _08477_/Y _08599_/A VGND VGND VPWR VPWR _08587_/A sky130_fd_sc_hd__o22a_1
XFILLER_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09108_ _09539_/B _09030_/B _09031_/B VGND VGND VPWR VPWR _09108_/Y sky130_fd_sc_hd__a21boi_1
X_10380_ _11805_/A _10453_/B _10379_/Y VGND VGND VPWR VPWR _10381_/A sky130_fd_sc_hd__o21ai_2
X_09039_ _09529_/B _09038_/B _09155_/B VGND VGND VPWR VPWR _09040_/A sky130_fd_sc_hd__a21bo_1
XFILLER_117_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12050_ _12040_/Y _12048_/X _12049_/Y VGND VGND VPWR VPWR _12050_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11001_ _11002_/A _11003_/B VGND VGND VPWR VPWR _11004_/A sky130_fd_sc_hd__and2_1
XFILLER_77_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15740_ _15752_/A _15740_/B VGND VGND VPWR VPWR _16110_/A sky130_fd_sc_hd__nor2_1
XFILLER_73_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12952_ _12952_/A _12951_/X VGND VGND VPWR VPWR _12952_/X sky130_fd_sc_hd__or2b_1
XFILLER_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15671_ _15671_/A _15671_/B VGND VGND VPWR VPWR _15671_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11903_ _11903_/A VGND VGND VPWR VPWR _11903_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14622_ _15341_/A _14656_/B VGND VGND VPWR VPWR _14622_/Y sky130_fd_sc_hd__nor2_1
X_12883_ _14532_/A _12938_/B VGND VGND VPWR VPWR _12883_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _13610_/A _11833_/B _10623_/A _11833_/Y VGND VGND VPWR VPWR _11834_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14553_ _14553_/A _14516_/X VGND VGND VPWR VPWR _14553_/X sky130_fd_sc_hd__or2b_1
XFILLER_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11765_ _11765_/A _11764_/X VGND VGND VPWR VPWR _11765_/X sky130_fd_sc_hd__or2b_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14484_ _15196_/A _14520_/B VGND VGND VPWR VPWR _14545_/A sky130_fd_sc_hd__and2_1
X_10716_ _11945_/A VGND VGND VPWR VPWR _13073_/A sky130_fd_sc_hd__buf_1
X_11696_ _11692_/Y _11695_/X _11692_/Y _11695_/X VGND VGND VPWR VPWR _11696_/X sky130_fd_sc_hd__a2bb2o_1
X_13504_ _13504_/A _13504_/B VGND VGND VPWR VPWR _13504_/Y sky130_fd_sc_hd__nand2_1
X_16223_ _16223_/A VGND VGND VPWR VPWR _16223_/Y sky130_fd_sc_hd__inv_2
X_13435_ _13361_/X _13434_/X _13361_/X _13434_/X VGND VGND VPWR VPWR _13435_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10647_ _10647_/A VGND VGND VPWR VPWR _10647_/Y sky130_fd_sc_hd__inv_2
Xrebuffer4 _16238_/A VGND VGND VPWR VPWR _16247_/C1 sky130_fd_sc_hd__dlymetal6s2s_1
X_16154_ _16270_/A _16336_/A VGND VGND VPWR VPWR _16154_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13366_ _13388_/A _13364_/X _13365_/X VGND VGND VPWR VPWR _13366_/X sky130_fd_sc_hd__o21a_1
X_10578_ _10539_/X _10577_/X _10539_/X _10577_/X VGND VGND VPWR VPWR _10651_/B sky130_fd_sc_hd__a2bb2o_1
X_16085_ _16082_/Y _16233_/A _16084_/Y VGND VGND VPWR VPWR _16089_/B sky130_fd_sc_hd__o21ai_1
X_12317_ _12235_/X _12316_/Y _12235_/A _12316_/Y VGND VGND VPWR VPWR _12318_/B sky130_fd_sc_hd__a2bb2o_1
X_13297_ _14739_/A _13297_/B VGND VGND VPWR VPWR _13297_/Y sky130_fd_sc_hd__nand2_1
X_15105_ _15105_/A _15104_/X VGND VGND VPWR VPWR _15105_/X sky130_fd_sc_hd__or2b_1
XFILLER_114_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12248_ _12201_/A _12154_/X _12200_/X VGND VGND VPWR VPWR _12248_/X sky130_fd_sc_hd__o21a_1
X_15036_ _15036_/A _15036_/B VGND VGND VPWR VPWR _15036_/X sky130_fd_sc_hd__or2_1
XFILLER_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12179_ _12179_/A _12179_/B VGND VGND VPWR VPWR _12179_/X sky130_fd_sc_hd__or2_1
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15938_ _15889_/X _15937_/Y _15889_/X _15937_/Y VGND VGND VPWR VPWR _15952_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15869_ _15869_/A VGND VGND VPWR VPWR _15894_/A sky130_fd_sc_hd__inv_2
XFILLER_37_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08410_ _08409_/A _08354_/Y _08409_/Y _08354_/A _08419_/A VGND VGND VPWR VPWR _09225_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09390_ _09344_/X _09389_/X _09344_/X _09389_/X VGND VGND VPWR VPWR _10420_/B sky130_fd_sc_hd__a2bb2o_4
X_08341_ input30/X _08341_/B VGND VGND VPWR VPWR _08342_/B sky130_fd_sc_hd__nor2_1
X_08272_ _08272_/A input11/X VGND VGND VPWR VPWR _08364_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09726_ _09770_/A _09770_/B _09725_/Y VGND VGND VPWR VPWR _09727_/A sky130_fd_sc_hd__o21ai_1
XFILLER_55_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09657_ _09603_/Y _09655_/X _09656_/Y VGND VGND VPWR VPWR _09657_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08608_ _08716_/B VGND VGND VPWR VPWR _08610_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09588_ _09989_/A VGND VGND VPWR VPWR _09990_/A sky130_fd_sc_hd__buf_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08538_/A _08323_/Y _08538_/Y _08323_/A VGND VGND VPWR VPWR _08540_/B sky130_fd_sc_hd__o22a_1
XFILLER_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11550_ _13883_/A _11649_/B _11549_/Y VGND VGND VPWR VPWR _11550_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10501_ _10500_/A _10499_/Y _10500_/Y _10499_/A _09941_/A VGND VGND VPWR VPWR _12926_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13220_ _14771_/A _13303_/B VGND VGND VPWR VPWR _13220_/Y sky130_fd_sc_hd__nor2_1
X_11481_ _11480_/A _11480_/B _11480_/X _11277_/X VGND VGND VPWR VPWR _11481_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10432_ _12825_/A _10432_/B VGND VGND VPWR VPWR _10432_/X sky130_fd_sc_hd__or2_1
X_13151_ _15243_/A _13119_/B _13119_/Y VGND VGND VPWR VPWR _13151_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10363_ _09971_/A _10362_/Y _09971_/Y _10362_/A _10446_/A VGND VGND VPWR VPWR _11755_/A
+ sky130_fd_sc_hd__o221a_1
X_13082_ _15258_/A _13109_/B VGND VGND VPWR VPWR _13082_/Y sky130_fd_sc_hd__nor2_1
X_12102_ _13053_/A _12158_/B _12101_/Y VGND VGND VPWR VPWR _12102_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12033_ _11967_/X _12032_/Y _11967_/X _12032_/Y VGND VGND VPWR VPWR _12053_/B sky130_fd_sc_hd__a2bb2o_1
X_10294_ _10335_/B VGND VGND VPWR VPWR _10294_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15723_ _15685_/A _15685_/B _15685_/Y VGND VGND VPWR VPWR _15723_/Y sky130_fd_sc_hd__o21ai_1
X_13984_ _13985_/A _13985_/B VGND VGND VPWR VPWR _13986_/A sky130_fd_sc_hd__and2_1
X_12935_ _12891_/Y _12933_/X _12934_/Y VGND VGND VPWR VPWR _12935_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15654_ _15667_/A _15667_/B VGND VGND VPWR VPWR _15785_/A sky130_fd_sc_hd__and2_1
XFILLER_61_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12866_ _12859_/X _12865_/Y _12859_/X _12865_/Y VGND VGND VPWR VPWR _12947_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15585_ _15685_/A _15685_/B VGND VGND VPWR VPWR _15585_/Y sky130_fd_sc_hd__nor2_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14605_/A _14604_/X VGND VGND VPWR VPWR _14605_/X sky130_fd_sc_hd__or2b_1
X_11817_ _11797_/X _11816_/X _11797_/X _11816_/X VGND VGND VPWR VPWR _11843_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _15190_/A _14536_/B VGND VGND VPWR VPWR _14536_/X sky130_fd_sc_hd__or2_1
X_12797_ _12780_/X _12796_/Y _12780_/X _12796_/Y VGND VGND VPWR VPWR _12856_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11748_ _10310_/A _11747_/A _10310_/Y _11759_/B VGND VGND VPWR VPWR _11750_/B sky130_fd_sc_hd__o22a_1
X_11679_ _11648_/A _11650_/X _11647_/X VGND VGND VPWR VPWR _11679_/X sky130_fd_sc_hd__o21a_1
X_14467_ _14467_/A _14467_/B VGND VGND VPWR VPWR _14467_/Y sky130_fd_sc_hd__nand2_1
X_16206_ _16104_/A _15805_/B _15805_/Y VGND VGND VPWR VPWR _16208_/A sky130_fd_sc_hd__o21ai_1
X_14398_ _15970_/A _14401_/B VGND VGND VPWR VPWR _15687_/A sky130_fd_sc_hd__and2_1
X_13418_ _14096_/A _13421_/B VGND VGND VPWR VPWR _13418_/Y sky130_fd_sc_hd__nor2_1
X_16137_ _16136_/A _16136_/B _16136_/X VGND VGND VPWR VPWR _16137_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13349_ _13349_/A _13349_/B VGND VGND VPWR VPWR _13349_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16068_ _16044_/A _16044_/B _16044_/Y VGND VGND VPWR VPWR _16068_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15019_ _11765_/X _15000_/X _11765_/X _15000_/X VGND VGND VPWR VPWR _15034_/B sky130_fd_sc_hd__a2bb2o_1
X_08890_ _08978_/A _08978_/B VGND VGND VPWR VPWR _08890_/X sky130_fd_sc_hd__and2_1
XFILLER_96_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09511_ _09494_/A _09494_/B _09494_/Y _09510_/X VGND VGND VPWR VPWR _09511_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09442_ _09198_/X _09360_/X _09198_/X _09360_/X VGND VGND VPWR VPWR _09442_/X sky130_fd_sc_hd__o2bb2a_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09373_ _09356_/X _09372_/X _09356_/X _09372_/X VGND VGND VPWR VPWR _09374_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08324_ _08324_/A VGND VGND VPWR VPWR _08324_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08255_ input16/X VGND VGND VPWR VPWR _08331_/A sky130_fd_sc_hd__inv_2
XFILLER_118_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09709_ _09709_/A _09709_/B VGND VGND VPWR VPWR _09709_/Y sky130_fd_sc_hd__nand2_1
X_10981_ _10981_/A _10981_/B VGND VGND VPWR VPWR _10981_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12720_ _12682_/A _12682_/B _12682_/Y _12719_/X VGND VGND VPWR VPWR _12720_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12651_ _12641_/Y _12649_/Y _14163_/B VGND VGND VPWR VPWR _12651_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_90_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11602_ _09749_/X _10034_/B _10034_/Y VGND VGND VPWR VPWR _11602_/X sky130_fd_sc_hd__o21a_1
X_12582_ _12582_/A VGND VGND VPWR VPWR _12582_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15370_ _15344_/X _15369_/X _15344_/X _15369_/X VGND VGND VPWR VPWR _15412_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14321_ _14335_/A _14321_/B VGND VGND VPWR VPWR _15960_/A sky130_fd_sc_hd__or2_1
X_11533_ _11533_/A _11533_/B VGND VGND VPWR VPWR _11533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14252_ _14234_/Y _14250_/Y _14251_/Y VGND VGND VPWR VPWR _14253_/A sky130_fd_sc_hd__o21ai_2
X_11464_ _14144_/A VGND VGND VPWR VPWR _13448_/A sky130_fd_sc_hd__buf_1
XFILLER_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13203_ _13150_/Y _13201_/X _13202_/Y VGND VGND VPWR VPWR _13203_/X sky130_fd_sc_hd__o21a_1
X_10415_ _12825_/A _10432_/B VGND VGND VPWR VPWR _10512_/A sky130_fd_sc_hd__and2_1
XFILLER_124_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14183_ _14282_/A _14183_/B VGND VGND VPWR VPWR _15857_/A sky130_fd_sc_hd__or2_1
XFILLER_109_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11395_ _11395_/A VGND VGND VPWR VPWR _11395_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13134_ _13967_/A VGND VGND VPWR VPWR _15167_/A sky130_fd_sc_hd__buf_1
X_10346_ _10903_/A _10346_/B VGND VGND VPWR VPWR _10347_/A sky130_fd_sc_hd__or2_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13065_/A _13024_/X VGND VGND VPWR VPWR _13065_/X sky130_fd_sc_hd__or2b_1
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ _10277_/A VGND VGND VPWR VPWR _10277_/Y sky130_fd_sc_hd__inv_2
X_12016_ _13063_/A _11976_/B _11976_/Y VGND VGND VPWR VPWR _12016_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13967_ _13967_/A _13968_/B VGND VGND VPWR VPWR _13969_/A sky130_fd_sc_hd__and2_1
X_15706_ _16125_/A _15823_/B VGND VGND VPWR VPWR _15706_/X sky130_fd_sc_hd__and2_1
X_12918_ _12835_/X _12915_/Y _12916_/Y _12917_/X VGND VGND VPWR VPWR _12920_/B sky130_fd_sc_hd__o22a_1
X_15637_ _14381_/X _15636_/X _14381_/X _15636_/X VGND VGND VPWR VPWR _15671_/B sky130_fd_sc_hd__a2bb2o_1
X_13898_ _13898_/A VGND VGND VPWR VPWR _15414_/A sky130_fd_sc_hd__buf_1
X_12849_ _12810_/Y _12847_/X _12848_/Y VGND VGND VPWR VPWR _12849_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _15562_/X _15567_/Y _15562_/X _15567_/Y VGND VGND VPWR VPWR _15568_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15499_ _15482_/X _15498_/X _15482_/X _15498_/X VGND VGND VPWR VPWR _15546_/B sky130_fd_sc_hd__a2bb2o_1
X_14519_ _14549_/A _14517_/X _14518_/X VGND VGND VPWR VPWR _14519_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09991_ _09967_/Y _09989_/Y _09990_/Y VGND VGND VPWR VPWR _09993_/B sky130_fd_sc_hd__o21ai_2
XFILLER_130_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08942_ _08942_/A _08942_/B VGND VGND VPWR VPWR _08942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08873_ _08762_/A _10133_/A _08762_/Y VGND VGND VPWR VPWR _08873_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09425_ _09266_/A _09423_/Y _09424_/Y VGND VGND VPWR VPWR _09433_/B sky130_fd_sc_hd__o21ai_1
XFILLER_40_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09356_ _08690_/A _09860_/A _09353_/Y _09355_/X VGND VGND VPWR VPWR _09356_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08307_ _08307_/A _08307_/B VGND VGND VPWR VPWR _08308_/A sky130_fd_sc_hd__or2_1
X_09287_ _09255_/Y _08954_/Y _09255_/Y _08954_/Y VGND VGND VPWR VPWR _10245_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08238_ _08238_/A _08238_/B VGND VGND VPWR VPWR _08239_/A sky130_fd_sc_hd__or2_1
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10200_ _10108_/A _10109_/A _10108_/Y _10109_/Y _10346_/B VGND VGND VPWR VPWR _10213_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11180_ _09436_/A _09141_/B _09141_/Y VGND VGND VPWR VPWR _11181_/A sky130_fd_sc_hd__o21ai_1
XFILLER_121_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10131_ _10131_/A _10131_/B VGND VGND VPWR VPWR _10132_/B sky130_fd_sc_hd__or2_1
XFILLER_125_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10062_ _10020_/X _10061_/Y _10020_/X _10061_/Y VGND VGND VPWR VPWR _10063_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14870_ _14825_/X _14869_/X _14825_/X _14869_/X VGND VGND VPWR VPWR _14924_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13821_ _14627_/A _13846_/B VGND VGND VPWR VPWR _13821_/Y sky130_fd_sc_hd__nor2_1
X_13752_ _11959_/X _13751_/X _11959_/X _13751_/X VGND VGND VPWR VPWR _13753_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12703_ _12703_/A _12703_/B VGND VGND VPWR VPWR _12703_/X sky130_fd_sc_hd__and2_1
X_10964_ _12082_/A _10964_/B VGND VGND VPWR VPWR _10964_/Y sky130_fd_sc_hd__nor2_1
X_16471_ _08229_/A _16471_/D VGND VGND VPWR VPWR _16471_/Q sky130_fd_sc_hd__dfxtp_1
X_10895_ _12049_/A VGND VGND VPWR VPWR _13829_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13683_ _13002_/X _13682_/X _13002_/A _13682_/X VGND VGND VPWR VPWR _13684_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12634_ _14184_/A _12632_/X _12633_/X VGND VGND VPWR VPWR _12634_/X sky130_fd_sc_hd__o21a_1
X_15422_ _15422_/A _15422_/B VGND VGND VPWR VPWR _15422_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12565_ _15529_/A VGND VGND VPWR VPWR _14912_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15353_ _15353_/A _15353_/B VGND VGND VPWR VPWR _15353_/X sky130_fd_sc_hd__or2_1
XFILLER_129_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14304_ _15906_/A _14278_/B _14278_/Y VGND VGND VPWR VPWR _14304_/Y sky130_fd_sc_hd__o21ai_1
X_11516_ _11516_/A _12273_/A VGND VGND VPWR VPWR _11516_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12496_ _12489_/X _12495_/X _12489_/X _12495_/X VGND VGND VPWR VPWR _12496_/X sky130_fd_sc_hd__a2bb2o_1
X_15284_ _14953_/A _15234_/B _15234_/Y _15283_/X VGND VGND VPWR VPWR _15284_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_8_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14235_ _14235_/A _14235_/B VGND VGND VPWR VPWR _15839_/A sky130_fd_sc_hd__nor2_1
X_11447_ _11442_/Y _12554_/A _11446_/Y VGND VGND VPWR VPWR _11453_/B sky130_fd_sc_hd__o21ai_1
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14166_ _15974_/A _14166_/B VGND VGND VPWR VPWR _14166_/X sky130_fd_sc_hd__or2_1
XFILLER_98_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11378_ _08901_/X _11378_/B VGND VGND VPWR VPWR _11378_/X sky130_fd_sc_hd__and2b_1
XFILLER_124_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13117_ _15246_/A _13117_/B VGND VGND VPWR VPWR _13117_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _09955_/A _09955_/B _09955_/X VGND VGND VPWR VPWR _10330_/A sky130_fd_sc_hd__o21ba_1
X_14097_ _14093_/Y _14095_/Y _14096_/Y VGND VGND VPWR VPWR _14101_/B sky130_fd_sc_hd__o21ai_2
XFILLER_79_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13048_ _13048_/A VGND VGND VPWR VPWR _13775_/A sky130_fd_sc_hd__inv_2
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14999_ _12703_/A _11743_/Y _11736_/Y _14998_/X VGND VGND VPWR VPWR _14999_/X sky130_fd_sc_hd__o22a_1
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09210_ _09857_/A VGND VGND VPWR VPWR _09731_/A sky130_fd_sc_hd__inv_2
X_09141_ _09436_/A _09141_/B VGND VGND VPWR VPWR _09141_/Y sky130_fd_sc_hd__nand2_1
X_09072_ _10017_/B _09072_/B VGND VGND VPWR VPWR _09073_/B sky130_fd_sc_hd__or2_1
XFILLER_30_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09974_ _09974_/A _09975_/B VGND VGND VPWR VPWR _09974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08925_ _08930_/A _09541_/A VGND VGND VPWR VPWR _09817_/A sky130_fd_sc_hd__or2_1
XFILLER_85_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08856_ _08934_/A _08856_/B VGND VGND VPWR VPWR _09460_/A sky130_fd_sc_hd__or2_1
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08787_ _09324_/A VGND VGND VPWR VPWR _09490_/A sky130_fd_sc_hd__buf_1
XFILLER_72_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10680_ _10680_/A VGND VGND VPWR VPWR _10680_/Y sky130_fd_sc_hd__inv_2
X_09408_ _09297_/A _10892_/A _09407_/X VGND VGND VPWR VPWR _09409_/B sky130_fd_sc_hd__o21ai_1
X_09339_ _09448_/A _09339_/B VGND VGND VPWR VPWR _09339_/X sky130_fd_sc_hd__or2_1
XFILLER_126_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12350_ _12346_/Y _12549_/A _12349_/Y VGND VGND VPWR VPWR _12541_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11301_ _12365_/A VGND VGND VPWR VPWR _13789_/A sky130_fd_sc_hd__buf_1
X_12281_ _13789_/A _12365_/B VGND VGND VPWR VPWR _12281_/Y sky130_fd_sc_hd__nand2_1
X_11232_ _14809_/A VGND VGND VPWR VPWR _12227_/A sky130_fd_sc_hd__inv_2
X_14020_ _13951_/X _14019_/Y _13951_/X _14019_/Y VGND VGND VPWR VPWR _14056_/B sky130_fd_sc_hd__a2bb2o_1
X_11163_ _11129_/X _11162_/X _11129_/X _11162_/X VGND VGND VPWR VPWR _11295_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10114_ _10114_/A _10114_/B VGND VGND VPWR VPWR _10115_/A sky130_fd_sc_hd__or2_1
XFILLER_121_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15971_ _15918_/Y _15969_/Y _15970_/Y VGND VGND VPWR VPWR _15971_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11094_ _11186_/A _11092_/X _11093_/X VGND VGND VPWR VPWR _11094_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14922_ _15546_/A _14922_/B VGND VGND VPWR VPWR _14922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10045_ _10026_/X _10044_/Y _10026_/X _10044_/Y VGND VGND VPWR VPWR _10081_/B sky130_fd_sc_hd__a2bb2o_1
X_14853_ _14834_/X _14852_/Y _14834_/X _14852_/Y VGND VGND VPWR VPWR _14958_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13804_ _13804_/A _13773_/X VGND VGND VPWR VPWR _13804_/X sky130_fd_sc_hd__or2b_1
XFILLER_36_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14784_ _14784_/A _14737_/X VGND VGND VPWR VPWR _14784_/X sky130_fd_sc_hd__or2b_1
XFILLER_44_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11996_ _11997_/A _11997_/B VGND VGND VPWR VPWR _11998_/A sky130_fd_sc_hd__and2_1
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13735_ _13767_/A _13767_/B VGND VGND VPWR VPWR _13813_/A sky130_fd_sc_hd__and2_1
XFILLER_44_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10947_ _10947_/A _10947_/B VGND VGND VPWR VPWR _10947_/Y sky130_fd_sc_hd__nor2_1
X_16454_ _16454_/A _16454_/B _16404_/B VGND VGND VPWR VPWR _16454_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_71_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13666_ _13628_/A _13665_/Y _13628_/A _13665_/Y VGND VGND VPWR VPWR _13695_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12617_ _12617_/A _12617_/B VGND VGND VPWR VPWR _14232_/B sky130_fd_sc_hd__or2_1
X_15405_ _15459_/A _15403_/X _15404_/X VGND VGND VPWR VPWR _15405_/X sky130_fd_sc_hd__o21a_1
X_10878_ _09286_/Y _10877_/A _09286_/A _10877_/Y _09445_/A VGND VGND VPWR VPWR _12053_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16385_ _16136_/A _16136_/B _16136_/X _16274_/Y VGND VGND VPWR VPWR _16385_/X sky130_fd_sc_hd__a22o_1
X_13597_ _13560_/A _13560_/B _13561_/A VGND VGND VPWR VPWR _13597_/Y sky130_fd_sc_hd__o21ai_1
X_12548_ _12544_/Y _12547_/Y _12544_/A _12547_/A _11707_/A VGND VGND VPWR VPWR _12627_/A
+ sky130_fd_sc_hd__o221a_1
X_15336_ _15384_/A _15334_/X _15335_/X VGND VGND VPWR VPWR _15336_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12479_ _12476_/Y _12477_/Y _12478_/Y VGND VGND VPWR VPWR _12479_/Y sky130_fd_sc_hd__o21ai_1
X_15267_ _15272_/A _15272_/B VGND VGND VPWR VPWR _15324_/A sky130_fd_sc_hd__and2_1
XANTENNA_2 input31/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14218_ _14095_/Y _14217_/X _14095_/Y _14217_/X VGND VGND VPWR VPWR _14219_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15198_ _15151_/X _15197_/Y _15151_/X _15197_/Y VGND VGND VPWR VPWR _15199_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14149_ _14149_/A _14149_/B VGND VGND VPWR VPWR _14149_/Y sky130_fd_sc_hd__nor2_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _08710_/A _09474_/B VGND VGND VPWR VPWR _08710_/Y sky130_fd_sc_hd__nor2_1
X_09690_ _09690_/A _09690_/B VGND VGND VPWR VPWR _09693_/B sky130_fd_sc_hd__or2_1
XFILLER_67_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08641_ _08719_/B VGND VGND VPWR VPWR _09230_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer25 _10191_/X VGND VGND VPWR VPWR _11525_/B1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer14 rebuffer15/X VGND VGND VPWR VPWR rebuffer14/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_35_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08572_ _08572_/A _10116_/B VGND VGND VPWR VPWR _08573_/A sky130_fd_sc_hd__or2_1
XFILLER_35_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09124_ _09120_/Y _09122_/Y _09123_/Y VGND VGND VPWR VPWR _09126_/B sky130_fd_sc_hd__o21ai_1
XFILLER_108_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09055_ _08773_/Y _09054_/A _08773_/A _09054_/Y VGND VGND VPWR VPWR _10011_/B sky130_fd_sc_hd__o22a_1
XFILLER_116_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09957_ _09957_/A _09958_/B VGND VGND VPWR VPWR _09957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08908_ _09549_/A _08609_/A _08611_/A VGND VGND VPWR VPWR _08908_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09888_/A _09888_/B VGND VGND VPWR VPWR _09888_/X sky130_fd_sc_hd__or2_1
XFILLER_73_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08839_ _08839_/A VGND VGND VPWR VPWR _08839_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11850_ _11850_/A VGND VGND VPWR VPWR _11913_/A sky130_fd_sc_hd__inv_2
X_11781_ _12825_/A VGND VGND VPWR VPWR _11787_/A sky130_fd_sc_hd__inv_2
X_10801_ _11916_/A _10801_/B VGND VGND VPWR VPWR _10801_/X sky130_fd_sc_hd__and2_1
XFILLER_26_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13520_ _13522_/A VGND VGND VPWR VPWR _15034_/A sky130_fd_sc_hd__buf_1
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10732_ _10732_/A VGND VGND VPWR VPWR _10732_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13451_ _13375_/Y _13449_/X _13450_/Y VGND VGND VPWR VPWR _13451_/X sky130_fd_sc_hd__o21a_1
X_10663_ _11850_/A _10663_/B VGND VGND VPWR VPWR _10663_/X sky130_fd_sc_hd__and2_1
X_16170_ _16266_/A _16332_/A VGND VGND VPWR VPWR _16170_/Y sky130_fd_sc_hd__nor2_1
X_13382_ _13382_/A _13369_/X VGND VGND VPWR VPWR _13382_/X sky130_fd_sc_hd__or2b_1
X_12402_ _12402_/A _12401_/X VGND VGND VPWR VPWR _12402_/X sky130_fd_sc_hd__or2b_1
X_10594_ _11901_/A _10638_/B VGND VGND VPWR VPWR _10594_/Y sky130_fd_sc_hd__nor2_1
X_12333_ _12239_/X _12332_/Y _12239_/X _12332_/Y VGND VGND VPWR VPWR _12580_/A sky130_fd_sc_hd__a2bb2o_1
X_15121_ _15095_/X _15120_/Y _15095_/X _15120_/Y VGND VGND VPWR VPWR _15122_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15052_ _15052_/A _15051_/X VGND VGND VPWR VPWR _15052_/X sky130_fd_sc_hd__or2b_1
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14003_ _14068_/A _14068_/B VGND VGND VPWR VPWR _14147_/A sky130_fd_sc_hd__and2_1
X_12264_ _13501_/A VGND VGND VPWR VPWR _12369_/A sky130_fd_sc_hd__inv_2
XFILLER_5_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11215_ _12218_/A VGND VGND VPWR VPWR _14028_/A sky130_fd_sc_hd__buf_1
X_12195_ _12159_/X _12194_/Y _12159_/X _12194_/Y VGND VGND VPWR VPWR _12249_/B sky130_fd_sc_hd__a2bb2o_1
X_11146_ _10240_/B _10147_/B _10147_/Y VGND VGND VPWR VPWR _11147_/A sky130_fd_sc_hd__a21oi_1
X_15954_ _15954_/A _15954_/B VGND VGND VPWR VPWR _15954_/X sky130_fd_sc_hd__or2_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11077_ _11240_/A _11074_/X _11076_/X VGND VGND VPWR VPWR _11077_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14905_ _14904_/A _14904_/B _12610_/A _14904_/Y VGND VGND VPWR VPWR _14905_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10028_ _09333_/A _08778_/B _10041_/B _10027_/X VGND VGND VPWR VPWR _10028_/X sky130_fd_sc_hd__o22a_1
X_15885_ _15885_/A _15885_/B VGND VGND VPWR VPWR _15885_/X sky130_fd_sc_hd__or2_1
XFILLER_91_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14836_ _14836_/A VGND VGND VPWR VPWR _15178_/A sky130_fd_sc_hd__buf_1
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14767_ _15351_/A _14830_/B VGND VGND VPWR VPWR _14767_/Y sky130_fd_sc_hd__nand2_1
X_11979_ _11979_/A VGND VGND VPWR VPWR _11979_/Y sky130_fd_sc_hd__inv_2
X_13718_ _13778_/A _13717_/Y _13778_/A _13717_/Y VGND VGND VPWR VPWR _13720_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14698_ _14657_/X _14697_/Y _14657_/X _14697_/Y VGND VGND VPWR VPWR _14735_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16437_ _16467_/Q _16437_/B _16465_/Q _16437_/D VGND VGND VPWR VPWR _16437_/X sky130_fd_sc_hd__or4_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13649_ _13649_/A _13649_/B VGND VGND VPWR VPWR _13709_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16368_ _16357_/X _16463_/Q _16358_/X _16407_/A _16361_/X VGND VGND VPWR VPWR _16463_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15319_ _15274_/X _15318_/Y _15274_/X _15318_/Y VGND VGND VPWR VPWR _15335_/B sky130_fd_sc_hd__a2bb2o_1
X_16299_ _16326_/A _16326_/B VGND VGND VPWR VPWR _16299_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09811_ _08962_/X _08623_/A _09457_/Y _09810_/X VGND VGND VPWR VPWR _09811_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09742_ _09742_/A _09742_/B VGND VGND VPWR VPWR _09745_/A sky130_fd_sc_hd__or2_1
XFILLER_101_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09673_ _09984_/A _09656_/B _09656_/Y VGND VGND VPWR VPWR _09673_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08624_ _08624_/A VGND VGND VPWR VPWR _08624_/Y sky130_fd_sc_hd__inv_2
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08555_ _10011_/A _08555_/B VGND VGND VPWR VPWR _09859_/A sky130_fd_sc_hd__or2_2
XFILLER_35_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08486_ _08269_/A _08352_/B _08478_/Y _08612_/A VGND VGND VPWR VPWR _08599_/A sky130_fd_sc_hd__o22a_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09107_ _09714_/A _09107_/B VGND VGND VPWR VPWR _09107_/X sky130_fd_sc_hd__and2_1
XFILLER_108_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09038_ _09529_/B _09038_/B VGND VGND VPWR VPWR _09155_/B sky130_fd_sc_hd__or2_1
X_11000_ _10929_/X _10999_/Y _10929_/X _10999_/Y VGND VGND VPWR VPWR _11003_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12951_ _14948_/A _12951_/B VGND VGND VPWR VPWR _12951_/X sky130_fd_sc_hd__or2_1
XFILLER_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15670_ _15646_/Y _15668_/Y _15669_/Y VGND VGND VPWR VPWR _15670_/X sky130_fd_sc_hd__o21a_1
X_11902_ _11876_/Y _11900_/Y _11901_/Y VGND VGND VPWR VPWR _11903_/A sky130_fd_sc_hd__o21ai_1
X_12882_ _12851_/X _12881_/Y _12851_/X _12881_/Y VGND VGND VPWR VPWR _12938_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14621_ _14583_/X _14620_/Y _14583_/X _14620_/Y VGND VGND VPWR VPWR _14656_/B sky130_fd_sc_hd__a2bb2o_1
X_11833_ _11833_/A _11833_/B VGND VGND VPWR VPWR _11833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _15258_/A VGND VGND VPWR VPWR _14580_/A sky130_fd_sc_hd__buf_1
XFILLER_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11764_ _11764_/A _11764_/B VGND VGND VPWR VPWR _11764_/X sky130_fd_sc_hd__or2_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _14468_/X _14482_/Y _14468_/X _14482_/Y VGND VGND VPWR VPWR _14520_/B sky130_fd_sc_hd__a2bb2o_1
X_11695_ _13463_/A _11629_/B _11629_/Y _11633_/X VGND VGND VPWR VPWR _11695_/X sky130_fd_sc_hd__o2bb2a_1
X_13503_ _11158_/X _13490_/X _11158_/X _13490_/X VGND VGND VPWR VPWR _13504_/B sky130_fd_sc_hd__o2bb2a_1
X_10715_ _10930_/A _10715_/B VGND VGND VPWR VPWR _11945_/A sky130_fd_sc_hd__or2_2
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16222_ _16089_/A _16089_/B _16089_/Y VGND VGND VPWR VPWR _16224_/A sky130_fd_sc_hd__o21ai_1
X_13434_ _13331_/A _13331_/B _13331_/A _13331_/B VGND VGND VPWR VPWR _13434_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10646_ _09773_/A _09773_/B _09773_/Y VGND VGND VPWR VPWR _10647_/A sky130_fd_sc_hd__o21ai_1
X_16153_ _16270_/B VGND VGND VPWR VPWR _16336_/A sky130_fd_sc_hd__buf_1
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer5 rebuffer6/X VGND VGND VPWR VPWR rebuffer5/X sky130_fd_sc_hd__dlygate4sd1_1
X_13365_ _13365_/A _13365_/B VGND VGND VPWR VPWR _13365_/X sky130_fd_sc_hd__or2_1
X_10577_ _10543_/X _10657_/B _10543_/X _10657_/B VGND VGND VPWR VPWR _10577_/X sky130_fd_sc_hd__a2bb2o_1
X_15104_ _15104_/A _15104_/B VGND VGND VPWR VPWR _15104_/X sky130_fd_sc_hd__or2_1
XFILLER_127_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16084_ _16084_/A _16084_/B VGND VGND VPWR VPWR _16084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12316_ _13351_/A _12236_/B _12236_/Y VGND VGND VPWR VPWR _12316_/Y sky130_fd_sc_hd__o21ai_1
X_13296_ _13296_/A VGND VGND VPWR VPWR _13296_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12247_ _14062_/A _12203_/B _12203_/Y _12246_/X VGND VGND VPWR VPWR _12247_/X sky130_fd_sc_hd__a2bb2o_1
X_15035_ _15073_/A _15033_/X _15034_/X VGND VGND VPWR VPWR _15035_/X sky130_fd_sc_hd__o21a_1
XFILLER_122_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12178_ _12179_/A _12179_/B VGND VGND VPWR VPWR _12180_/A sky130_fd_sc_hd__and2_1
XFILLER_122_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11129_ _11128_/A _11128_/B _11128_/X _10952_/X VGND VGND VPWR VPWR _11129_/X sky130_fd_sc_hd__o22a_1
X_15937_ _15890_/A _15890_/B _15890_/Y VGND VGND VPWR VPWR _15937_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15868_ _15896_/A _15896_/B VGND VGND VPWR VPWR _15868_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14819_ _14806_/A _14806_/B _14806_/X _14818_/X VGND VGND VPWR VPWR _14819_/X sky130_fd_sc_hd__o22a_1
XFILLER_91_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15799_ _15799_/A VGND VGND VPWR VPWR _16099_/A sky130_fd_sc_hd__buf_1
X_08340_ _08338_/Y _08339_/A _08338_/A _08339_/Y _08304_/A VGND VGND VPWR VPWR _09213_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08271_ input27/X VGND VGND VPWR VPWR _08272_/A sky130_fd_sc_hd__inv_2
XFILLER_32_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09725_ _09770_/A _09770_/B VGND VGND VPWR VPWR _09725_/Y sky130_fd_sc_hd__nand2_1
X_09656_ _09984_/A _09656_/B VGND VGND VPWR VPWR _09656_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08607_ _09456_/B VGND VGND VPWR VPWR _08716_/B sky130_fd_sc_hd__inv_2
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09587_ _09513_/X _09586_/X _09513_/X _09586_/X VGND VGND VPWR VPWR _09989_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08538_/A VGND VGND VPWR VPWR _08538_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08469_ input22/X input6/X VGND VGND VPWR VPWR _08469_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10500_ _10500_/A VGND VGND VPWR VPWR _10500_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11480_ _11480_/A _11480_/B VGND VGND VPWR VPWR _11480_/X sky130_fd_sc_hd__and2_1
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10431_ _12826_/A _10430_/B _10428_/X _10430_/X VGND VGND VPWR VPWR _10431_/X sky130_fd_sc_hd__o22a_1
XFILLER_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13150_ _13202_/A _13202_/B VGND VGND VPWR VPWR _13150_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10362_ _10362_/A VGND VGND VPWR VPWR _10362_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13081_ _13017_/X _13080_/X _13017_/X _13080_/X VGND VGND VPWR VPWR _13109_/B sky130_fd_sc_hd__a2bb2o_1
X_12101_ _12158_/A _12158_/B VGND VGND VPWR VPWR _12101_/Y sky130_fd_sc_hd__nand2_1
X_10293_ _10212_/X _12704_/A _10212_/X _12704_/A VGND VGND VPWR VPWR _10335_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12032_ _13083_/A _11968_/B _11968_/Y VGND VGND VPWR VPWR _12032_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13983_ _13980_/X _13982_/X _13980_/X _13982_/X VGND VGND VPWR VPWR _13985_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15722_ _16119_/A VGND VGND VPWR VPWR _15817_/A sky130_fd_sc_hd__inv_2
X_12934_ _12934_/A _12934_/B VGND VGND VPWR VPWR _12934_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15653_ _16030_/A VGND VGND VPWR VPWR _15667_/B sky130_fd_sc_hd__inv_2
XFILLER_73_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12865_ _13873_/A _12860_/B _12860_/Y VGND VGND VPWR VPWR _12865_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15584_ _14395_/X _15583_/X _14395_/X _15583_/X VGND VGND VPWR VPWR _15685_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _15187_/A _14604_/B VGND VGND VPWR VPWR _14604_/X sky130_fd_sc_hd__or2_1
X_11816_ _10441_/X _11845_/B _10441_/X _11845_/B VGND VGND VPWR VPWR _11816_/X sky130_fd_sc_hd__a2bb2o_1
X_12796_ _12781_/A _12781_/B _12781_/Y VGND VGND VPWR VPWR _12796_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _15190_/A _14536_/B VGND VGND VPWR VPWR _14537_/A sky130_fd_sc_hd__and2_1
X_11747_ _11747_/A VGND VGND VPWR VPWR _11759_/B sky130_fd_sc_hd__inv_2
X_16205_ _16205_/A _16205_/B VGND VGND VPWR VPWR _16255_/A sky130_fd_sc_hd__or2_1
X_11678_ _11655_/A _11580_/X _11654_/X VGND VGND VPWR VPWR _11678_/Y sky130_fd_sc_hd__o21ai_1
X_14466_ _14448_/Y _14464_/X _14465_/Y VGND VGND VPWR VPWR _14466_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14397_ _15583_/A _14395_/X _14396_/X VGND VGND VPWR VPWR _14401_/B sky130_fd_sc_hd__o21ai_1
X_13417_ _13413_/X _13415_/Y _14351_/B VGND VGND VPWR VPWR _13421_/B sky130_fd_sc_hd__o21ai_2
X_10629_ _11892_/A _10629_/B VGND VGND VPWR VPWR _10629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16136_ _16136_/A _16136_/B VGND VGND VPWR VPWR _16136_/X sky130_fd_sc_hd__or2_1
X_13348_ _13273_/X _13347_/Y _13273_/X _13347_/Y VGND VGND VPWR VPWR _13349_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16067_ _16114_/A _16114_/B VGND VGND VPWR VPWR _16067_/X sky130_fd_sc_hd__and2_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13279_ _14727_/A _13279_/B VGND VGND VPWR VPWR _13279_/Y sky130_fd_sc_hd__nand2_1
X_15018_ _15036_/A _15036_/B VGND VGND VPWR VPWR _15070_/A sky130_fd_sc_hd__and2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09510_ _09496_/A _09496_/B _09496_/Y _09509_/X VGND VGND VPWR VPWR _09510_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09441_ _09429_/A _09429_/B _09429_/X _09440_/X VGND VGND VPWR VPWR _09441_/X sky130_fd_sc_hd__a22o_2
X_09372_ _09474_/B _09861_/A _09351_/A VGND VGND VPWR VPWR _09372_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08323_ _08323_/A VGND VGND VPWR VPWR _08323_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08254_ input17/X _08254_/B VGND VGND VPWR VPWR _08327_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09708_ _09681_/A _09101_/A _08928_/A _09707_/Y VGND VGND VPWR VPWR _09709_/B sky130_fd_sc_hd__o22a_1
XFILLER_28_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10980_ _09328_/B _10241_/B _10241_/X VGND VGND VPWR VPWR _10981_/B sky130_fd_sc_hd__a21boi_1
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09639_ _09543_/X _09638_/Y _09543_/X _09638_/Y VGND VGND VPWR VPWR _10740_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12650_ _12650_/A _12650_/B VGND VGND VPWR VPWR _14163_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11601_ _11616_/A VGND VGND VPWR VPWR _12679_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14320_ _13437_/X _14319_/X _13437_/X _14319_/X VGND VGND VPWR VPWR _14321_/B sky130_fd_sc_hd__a2bb2oi_1
X_12581_ _14910_/A _12334_/B _12334_/Y VGND VGND VPWR VPWR _12582_/A sky130_fd_sc_hd__o21ai_1
XFILLER_128_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11532_ _09371_/B _10238_/B _10238_/X VGND VGND VPWR VPWR _11533_/B sky130_fd_sc_hd__a21boi_1
X_14251_ _15881_/A _14251_/B VGND VGND VPWR VPWR _14251_/Y sky130_fd_sc_hd__nand2_1
X_11463_ _12407_/A VGND VGND VPWR VPWR _14144_/A sky130_fd_sc_hd__buf_1
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14182_ _14122_/X _14181_/Y _14122_/X _14181_/Y VGND VGND VPWR VPWR _14183_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ _13202_/A _13202_/B VGND VGND VPWR VPWR _13202_/Y sky130_fd_sc_hd__nand2_1
X_10414_ _10357_/X _10413_/X _10357_/X _10413_/X VGND VGND VPWR VPWR _10432_/B sky130_fd_sc_hd__a2bb2o_1
X_13133_ _13133_/A VGND VGND VPWR VPWR _13967_/A sky130_fd_sc_hd__inv_2
XFILLER_3_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11394_ _08968_/A _08968_/B _08968_/Y VGND VGND VPWR VPWR _11395_/A sky130_fd_sc_hd__o21ai_1
XFILLER_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10345_ _10421_/A VGND VGND VPWR VPWR _10424_/A sky130_fd_sc_hd__inv_2
X_13064_ _13769_/A VGND VGND VPWR VPWR _15249_/A sky130_fd_sc_hd__buf_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10276_ _10228_/A _10228_/B _10228_/Y VGND VGND VPWR VPWR _10277_/A sky130_fd_sc_hd__a21oi_2
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ _12061_/A VGND VGND VPWR VPWR _13196_/A sky130_fd_sc_hd__buf_1
XFILLER_120_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13966_ _13543_/X _13965_/X _13543_/X _13965_/X VGND VGND VPWR VPWR _13968_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15705_ _15697_/X _15704_/Y _15697_/X _15704_/Y VGND VGND VPWR VPWR _15823_/B sky130_fd_sc_hd__a2bb2o_1
X_13897_ _15416_/A _13958_/B VGND VGND VPWR VPWR _13897_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12917_ _12836_/A _12836_/B _12836_/X VGND VGND VPWR VPWR _12917_/X sky130_fd_sc_hd__o21ba_1
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15636_ _15636_/A _14382_/X VGND VGND VPWR VPWR _15636_/X sky130_fd_sc_hd__or2b_1
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12848_ _12848_/A _12848_/B VGND VGND VPWR VPWR _12848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ _15565_/X _15566_/X _15565_/X _15566_/X VGND VGND VPWR VPWR _15567_/Y sky130_fd_sc_hd__a2bb2oi_1
X_12779_ _12779_/A _12779_/B VGND VGND VPWR VPWR _12779_/Y sky130_fd_sc_hd__nand2_1
X_15498_ _15446_/A _15446_/B _15446_/A _15446_/B VGND VGND VPWR VPWR _15498_/X sky130_fd_sc_hd__a2bb2o_1
X_14518_ _15199_/A _14518_/B VGND VGND VPWR VPWR _14518_/X sky130_fd_sc_hd__or2_1
X_14449_ _14425_/A _14425_/B _14425_/Y VGND VGND VPWR VPWR _14449_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16119_ _16119_/A _16119_/B VGND VGND VPWR VPWR _16119_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09990_ _09990_/A _09990_/B VGND VGND VPWR VPWR _09990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08941_ _08678_/A _08940_/X _08678_/A _08940_/X VGND VGND VPWR VPWR _11405_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08872_ _08693_/X _08871_/Y _08693_/X _08871_/Y VGND VGND VPWR VPWR _08984_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09424_ _09424_/A _09424_/B VGND VGND VPWR VPWR _09424_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09355_ _08688_/A _09859_/A _09354_/Y _09319_/X VGND VGND VPWR VPWR _09355_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09286_ _09286_/A VGND VGND VPWR VPWR _09286_/Y sky130_fd_sc_hd__inv_2
X_08306_ input22/X _08306_/B VGND VGND VPWR VPWR _08307_/B sky130_fd_sc_hd__nor2_1
X_08237_ _08237_/A input23/X VGND VGND VPWR VPWR _08238_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10130_ _10130_/A _10130_/B VGND VGND VPWR VPWR _10131_/B sky130_fd_sc_hd__or2_1
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10061_ _10061_/A _10061_/B VGND VGND VPWR VPWR _10061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13820_ _13762_/X _13819_/X _13762_/X _13819_/X VGND VGND VPWR VPWR _13846_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13751_ _13684_/A _13684_/B _13684_/A _13684_/B VGND VGND VPWR VPWR _13751_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10963_ _10960_/Y _12690_/A _10810_/X _10962_/Y VGND VGND VPWR VPWR _10963_/X sky130_fd_sc_hd__o22a_1
X_16470_ _08229_/A _16470_/D VGND VGND VPWR VPWR _16470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12702_ _10226_/X _12657_/Y _10226_/X _12657_/Y VGND VGND VPWR VPWR _12703_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15421_ _15435_/A _15419_/X _15420_/X VGND VGND VPWR VPWR _15421_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_70_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13682_ _13003_/A _13612_/A _13610_/Y _13612_/Y VGND VGND VPWR VPWR _13682_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10894_ _09297_/A _10893_/A _09297_/Y _10893_/Y _09445_/A VGND VGND VPWR VPWR _12049_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12633_ _12633_/A _12633_/B VGND VGND VPWR VPWR _12633_/X sky130_fd_sc_hd__or2_1
XFILLER_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12564_ _12564_/A VGND VGND VPWR VPWR _12564_/Y sky130_fd_sc_hd__inv_2
X_15352_ _15360_/A _15350_/X _15351_/X VGND VGND VPWR VPWR _15352_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14303_ _14309_/A _14303_/B VGND VGND VPWR VPWR _15966_/A sky130_fd_sc_hd__or2_1
X_15283_ _14833_/A _15237_/B _15237_/Y _15282_/X VGND VGND VPWR VPWR _15283_/X sky130_fd_sc_hd__a2bb2o_1
X_11515_ _12373_/A VGND VGND VPWR VPWR _12273_/A sky130_fd_sc_hd__inv_2
XFILLER_8_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14234_ _15881_/A _14251_/B VGND VGND VPWR VPWR _14234_/Y sky130_fd_sc_hd__nor2_1
X_12495_ _12492_/Y _12493_/Y _12494_/Y VGND VGND VPWR VPWR _12495_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11446_ _15534_/A _11446_/B VGND VGND VPWR VPWR _11446_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14165_ _15974_/A _14166_/B VGND VGND VPWR VPWR _14167_/A sky130_fd_sc_hd__and2_1
X_11377_ _12309_/A _11377_/B VGND VGND VPWR VPWR _11377_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14096_ _14096_/A _14096_/B VGND VGND VPWR VPWR _14096_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13116_ _13067_/Y _13114_/X _13115_/Y VGND VGND VPWR VPWR _13116_/X sky130_fd_sc_hd__o21a_1
X_10328_ _13528_/A _10328_/B VGND VGND VPWR VPWR _10328_/X sky130_fd_sc_hd__and2_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13047_ _14833_/A _13123_/B VGND VGND VPWR VPWR _13047_/Y sky130_fd_sc_hd__nor2_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10259_ _09263_/B _10242_/B _10242_/X _10826_/A VGND VGND VPWR VPWR _10981_/A sky130_fd_sc_hd__a22o_1
XFILLER_78_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14998_ _11731_/A _11730_/Y _11724_/Y _14997_/X VGND VGND VPWR VPWR _14998_/X sky130_fd_sc_hd__o22a_1
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13949_ _13917_/Y _13947_/X _13948_/Y VGND VGND VPWR VPWR _13949_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15619_ _16038_/A VGND VGND VPWR VPWR _15675_/A sky130_fd_sc_hd__inv_2
XFILLER_62_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09140_ _09140_/A VGND VGND VPWR VPWR _09140_/Y sky130_fd_sc_hd__inv_2
X_09071_ _10018_/B _09071_/B VGND VGND VPWR VPWR _09072_/B sky130_fd_sc_hd__or2_1
XFILLER_128_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09973_ _09963_/Y _09972_/Y _09960_/Y VGND VGND VPWR VPWR _09975_/B sky130_fd_sc_hd__o21ai_2
XFILLER_131_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08924_ _09541_/A _10098_/B _08678_/A VGND VGND VPWR VPWR _08932_/B sky130_fd_sc_hd__o21ai_1
XFILLER_85_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08855_ _09503_/A _09041_/B VGND VGND VPWR VPWR _08855_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08786_ _09470_/A _08786_/B VGND VGND VPWR VPWR _08786_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09407_ _09407_/A _09407_/B VGND VGND VPWR VPWR _09407_/X sky130_fd_sc_hd__or2_1
X_09338_ _08762_/A _08760_/Y _10035_/A _09337_/X VGND VGND VPWR VPWR _09338_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_40_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11300_ _12944_/A VGND VGND VPWR VPWR _12365_/A sky130_fd_sc_hd__inv_2
X_09269_ _09269_/A _09269_/B VGND VGND VPWR VPWR _09269_/X sky130_fd_sc_hd__or2_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12280_ _12260_/X _12279_/X _12260_/X _12279_/X VGND VGND VPWR VPWR _12365_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11231_ _11231_/A _11249_/B VGND VGND VPWR VPWR _14809_/A sky130_fd_sc_hd__or2_1
XFILLER_122_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11162_ _12259_/A _11302_/B _12259_/A _11302_/B VGND VGND VPWR VPWR _11162_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10113_ _10113_/A _10113_/B VGND VGND VPWR VPWR _10114_/A sky130_fd_sc_hd__or2_1
X_15970_ _15970_/A _15970_/B VGND VGND VPWR VPWR _15970_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11093_ _13898_/A _11093_/B VGND VGND VPWR VPWR _11093_/X sky130_fd_sc_hd__or2_1
XFILLER_76_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14921_ _14879_/Y _14919_/X _14920_/Y VGND VGND VPWR VPWR _14921_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10044_ _10044_/A _10044_/B VGND VGND VPWR VPWR _10044_/Y sky130_fd_sc_hd__nor2_1
X_14852_ _14953_/A _14953_/B _14851_/Y VGND VGND VPWR VPWR _14852_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13803_ _14664_/A _13858_/B VGND VGND VPWR VPWR _13803_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14783_ _15449_/A VGND VGND VPWR VPWR _14786_/A sky130_fd_sc_hd__buf_1
X_11995_ _10823_/A _11994_/A _10823_/Y _12082_/B VGND VGND VPWR VPWR _11997_/B sky130_fd_sc_hd__o22a_1
XFILLER_90_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13734_ _13696_/X _13733_/X _13696_/X _13733_/X VGND VGND VPWR VPWR _13767_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10946_ _10946_/A VGND VGND VPWR VPWR _10946_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16453_ _16349_/X _16406_/A _16409_/A VGND VGND VPWR VPWR _16454_/B sky130_fd_sc_hd__o21a_1
XFILLER_71_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13665_ _15131_/A _13630_/B _13630_/Y VGND VGND VPWR VPWR _13665_/Y sky130_fd_sc_hd__o21ai_1
X_10877_ _10877_/A VGND VGND VPWR VPWR _10877_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16384_ _16160_/A _16384_/B VGND VGND VPWR VPWR _16395_/A sky130_fd_sc_hd__nand2b_1
X_12616_ _12616_/A VGND VGND VPWR VPWR _14236_/A sky130_fd_sc_hd__inv_2
X_15404_ _15404_/A _15404_/B VGND VGND VPWR VPWR _15404_/X sky130_fd_sc_hd__or2_1
X_15335_ _15335_/A _15335_/B VGND VGND VPWR VPWR _15335_/X sky130_fd_sc_hd__or2_1
X_13596_ _13629_/A _13630_/B VGND VGND VPWR VPWR _13596_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12547_ _12547_/A VGND VGND VPWR VPWR _12547_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12478_ _13995_/A _12478_/B VGND VGND VPWR VPWR _12478_/Y sky130_fd_sc_hd__nand2_1
X_15266_ _15217_/X _15265_/Y _15217_/X _15265_/Y VGND VGND VPWR VPWR _15272_/B sky130_fd_sc_hd__a2bb2o_1
XANTENNA_3 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11429_ _15519_/A _11429_/B VGND VGND VPWR VPWR _11429_/X sky130_fd_sc_hd__or2_1
X_14217_ _14096_/A _14096_/B _14096_/Y VGND VGND VPWR VPWR _14217_/X sky130_fd_sc_hd__o21a_1
X_15197_ _15131_/A _15131_/B _15131_/Y VGND VGND VPWR VPWR _15197_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14148_ _14067_/X _14147_/X _14067_/X _14147_/X VGND VGND VPWR VPWR _14149_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ _14114_/A _14115_/A VGND VGND VPWR VPWR _14079_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08640_ _09459_/B VGND VGND VPWR VPWR _08719_/B sky130_fd_sc_hd__inv_2
Xrebuffer26 _16231_/B VGND VGND VPWR VPWR _16309_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_66_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer15 rebuffer16/X VGND VGND VPWR VPWR rebuffer15/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08571_ _08571_/A VGND VGND VPWR VPWR _10116_/B sky130_fd_sc_hd__inv_2
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09123_ _09703_/A _09123_/B VGND VGND VPWR VPWR _09123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09054_ _09054_/A VGND VGND VPWR VPWR _09054_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09956_ _09955_/A _09955_/B _09954_/Y _09955_/X VGND VGND VPWR VPWR _09958_/B sky130_fd_sc_hd__o22ai_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09887_/A _09887_/B VGND VGND VPWR VPWR _09888_/B sky130_fd_sc_hd__or2_1
X_08907_ _08972_/A _08972_/B VGND VGND VPWR VPWR _08907_/X sky130_fd_sc_hd__and2_1
XFILLER_106_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _08718_/A _09462_/B _08718_/Y VGND VGND VPWR VPWR _08839_/A sky130_fd_sc_hd__a21oi_2
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08769_ _10010_/A VGND VGND VPWR VPWR _08770_/A sky130_fd_sc_hd__buf_1
XFILLER_82_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11780_ _11780_/A _11780_/B VGND VGND VPWR VPWR _11780_/X sky130_fd_sc_hd__and2_1
X_10800_ _10951_/A VGND VGND VPWR VPWR _11007_/A sky130_fd_sc_hd__buf_1
XFILLER_41_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10731_ _10731_/A VGND VGND VPWR VPWR _10731_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13450_ _13450_/A _13450_/B VGND VGND VPWR VPWR _13450_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12401_ _13545_/A _12401_/B VGND VGND VPWR VPWR _12401_/X sky130_fd_sc_hd__or2_1
X_10662_ _10795_/A VGND VGND VPWR VPWR _11014_/A sky130_fd_sc_hd__buf_1
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13381_ _14138_/A _13446_/B VGND VGND VPWR VPWR _13381_/Y sky130_fd_sc_hd__nor2_1
X_10593_ _10530_/X _10592_/Y _10530_/X _10592_/Y VGND VGND VPWR VPWR _10638_/B sky130_fd_sc_hd__a2bb2o_1
X_12332_ _12224_/A _12224_/B _12224_/Y VGND VGND VPWR VPWR _12332_/Y sky130_fd_sc_hd__o21ai_1
X_15120_ _15063_/A _15063_/B _15063_/Y VGND VGND VPWR VPWR _15120_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12263_ _12261_/A _12261_/B _12261_/X _12262_/Y VGND VGND VPWR VPWR _12369_/B sky130_fd_sc_hd__a22o_1
X_15051_ _15051_/A _15051_/B VGND VGND VPWR VPWR _15051_/X sky130_fd_sc_hd__or2_1
XFILLER_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11214_ _13334_/A VGND VGND VPWR VPWR _12218_/A sky130_fd_sc_hd__inv_2
X_14002_ _13963_/X _14001_/Y _13963_/X _14001_/Y VGND VGND VPWR VPWR _14068_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12194_ _13048_/A _12252_/B _12193_/Y VGND VGND VPWR VPWR _12194_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11145_ _11145_/A VGND VGND VPWR VPWR _12268_/A sky130_fd_sc_hd__inv_2
X_15953_ _16017_/A _15951_/X _15952_/X VGND VGND VPWR VPWR _15953_/X sky130_fd_sc_hd__o21a_1
X_11076_ _15392_/A _11076_/B VGND VGND VPWR VPWR _11076_/X sky130_fd_sc_hd__or2_1
X_14904_ _14904_/A _14904_/B VGND VGND VPWR VPWR _14904_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10027_ _09452_/A _08786_/B _10044_/B _10026_/X VGND VGND VPWR VPWR _10027_/X sky130_fd_sc_hd__o22a_1
X_15884_ _14243_/A _15839_/B _14237_/A _14371_/X _14243_/B VGND VGND VPWR VPWR _15885_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14835_ _14748_/X _14762_/A _14761_/X VGND VGND VPWR VPWR _14835_/X sky130_fd_sc_hd__o21a_1
XFILLER_17_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14766_ _14747_/X _14765_/Y _14747_/X _14765_/Y VGND VGND VPWR VPWR _14830_/B sky130_fd_sc_hd__a2bb2o_1
X_11978_ _11978_/A _11978_/B VGND VGND VPWR VPWR _11978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10929_ _13058_/A _10842_/B _10842_/Y _10776_/X VGND VGND VPWR VPWR _10929_/X sky130_fd_sc_hd__a2bb2o_1
X_13717_ _15116_/A _13779_/B _13716_/Y VGND VGND VPWR VPWR _13717_/Y sky130_fd_sc_hd__o21ai_1
X_14697_ _15343_/A _14658_/B _14658_/Y VGND VGND VPWR VPWR _14697_/Y sky130_fd_sc_hd__o21ai_1
X_16436_ _16460_/Q _16459_/Q _16465_/Q _16435_/X _16437_/D VGND VGND VPWR VPWR _16436_/X
+ sky130_fd_sc_hd__o41a_1
X_13648_ _13539_/X _13647_/Y _13539_/X _13647_/Y VGND VGND VPWR VPWR _13649_/B sky130_fd_sc_hd__a2bb2o_1
X_16367_ _16325_/X _16366_/Y _16325_/X _16366_/Y VGND VGND VPWR VPWR _16407_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13579_ _12846_/A _13556_/B _13557_/Y _13578_/X VGND VGND VPWR VPWR _13579_/X sky130_fd_sc_hd__o22a_1
X_16298_ _16259_/X _16297_/Y _16259_/X _16297_/Y VGND VGND VPWR VPWR _16326_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15318_ _14578_/A _15261_/B _15261_/Y VGND VGND VPWR VPWR _15318_/Y sky130_fd_sc_hd__o21ai_1
X_15249_ _15249_/A _15249_/B VGND VGND VPWR VPWR _15249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09810_ _09458_/Y _09809_/X _09462_/X VGND VGND VPWR VPWR _09810_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09741_ _08535_/A _09743_/B _08535_/A _09743_/B VGND VGND VPWR VPWR _09742_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09672_ _09672_/A VGND VGND VPWR VPWR _10930_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08623_ _08623_/A _10112_/B VGND VGND VPWR VPWR _08624_/A sky130_fd_sc_hd__or2_1
XFILLER_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _08554_/A VGND VGND VPWR VPWR _10011_/A sky130_fd_sc_hd__buf_1
XFILLER_52_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08485_ _08272_/A _08363_/B _08479_/Y _08625_/A VGND VGND VPWR VPWR _08612_/A sky130_fd_sc_hd__o22a_1
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09106_ _09407_/A _09104_/B _09104_/X _09105_/X VGND VGND VPWR VPWR _09107_/B sky130_fd_sc_hd__o22a_1
XFILLER_108_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09037_ _09531_/B _09037_/B VGND VGND VPWR VPWR _09038_/B sky130_fd_sc_hd__or2_1
XFILLER_124_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09939_ _09935_/Y _09938_/X _09935_/Y _09938_/X VGND VGND VPWR VPWR _11592_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12950_ _14948_/A _12951_/B VGND VGND VPWR VPWR _12952_/A sky130_fd_sc_hd__and2_1
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11901_ _11901_/A _11901_/B VGND VGND VPWR VPWR _11901_/Y sky130_fd_sc_hd__nand2_1
X_12881_ _12852_/A _12852_/B _12852_/Y VGND VGND VPWR VPWR _12881_/Y sky130_fd_sc_hd__o21ai_1
X_14620_ _14584_/A _14584_/B _14584_/Y VGND VGND VPWR VPWR _14620_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11832_ _11792_/X _11831_/X _11792_/X _11831_/X VGND VGND VPWR VPWR _11833_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14582_/A _14582_/B VGND VGND VPWR VPWR _14551_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11764_/A _11764_/B VGND VGND VPWR VPWR _11765_/A sky130_fd_sc_hd__and2_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _13995_/A VGND VGND VPWR VPWR _13463_/A sky130_fd_sc_hd__clkbuf_2
X_14482_ _14469_/A _14469_/B _14469_/Y VGND VGND VPWR VPWR _14482_/Y sky130_fd_sc_hd__o21ai_1
X_13502_ _13504_/A VGND VGND VPWR VPWR _15046_/A sky130_fd_sc_hd__buf_1
XFILLER_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10714_ _09651_/X _10713_/X _09651_/X _10713_/X VGND VGND VPWR VPWR _10715_/B sky130_fd_sc_hd__a2bb2oi_1
X_16221_ _16253_/A _16320_/A VGND VGND VPWR VPWR _16221_/Y sky130_fd_sc_hd__nor2_1
X_13433_ _14112_/A _13436_/B VGND VGND VPWR VPWR _13433_/Y sky130_fd_sc_hd__nor2_1
X_10645_ _10582_/Y _10643_/Y _10644_/Y VGND VGND VPWR VPWR _10782_/A sky130_fd_sc_hd__o21ai_1
XFILLER_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16152_ _16160_/A _16152_/B VGND VGND VPWR VPWR _16270_/B sky130_fd_sc_hd__or2_1
X_13364_ _13391_/A _13362_/X _13363_/X VGND VGND VPWR VPWR _13364_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12315_ _13405_/A VGND VGND VPWR VPWR _14082_/A sky130_fd_sc_hd__inv_2
X_15103_ _15104_/A _15104_/B VGND VGND VPWR VPWR _15105_/A sky130_fd_sc_hd__and2_1
X_10576_ _10545_/X _10575_/X _10545_/X _10575_/X VGND VGND VPWR VPWR _10657_/B sky130_fd_sc_hd__a2bb2o_1
Xrebuffer6 rebuffer7/X VGND VGND VPWR VPWR rebuffer6/X sky130_fd_sc_hd__dlygate4sd1_1
X_16083_ _15778_/A _15765_/A _15781_/B VGND VGND VPWR VPWR _16233_/A sky130_fd_sc_hd__o21ai_2
X_13295_ _13235_/Y _13293_/Y _13294_/Y VGND VGND VPWR VPWR _13296_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12246_ _14060_/A _12206_/B _12206_/Y _12245_/X VGND VGND VPWR VPWR _12246_/X sky130_fd_sc_hd__a2bb2o_1
X_15034_ _15034_/A _15034_/B VGND VGND VPWR VPWR _15034_/X sky130_fd_sc_hd__or2_1
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12177_ _11152_/A _12176_/A _11152_/Y _12268_/B VGND VGND VPWR VPWR _12179_/B sky130_fd_sc_hd__o22a_1
XFILLER_110_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11128_ _11128_/A _11128_/B VGND VGND VPWR VPWR _11128_/X sky130_fd_sc_hd__and2_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15936_ _15954_/A _15954_/B VGND VGND VPWR VPWR _16014_/A sky130_fd_sc_hd__and2_1
X_11059_ _11792_/A VGND VGND VPWR VPWR _13936_/A sky130_fd_sc_hd__buf_1
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15867_ _14202_/X _15845_/X _14202_/X _15845_/X VGND VGND VPWR VPWR _15896_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14818_ _14809_/A _14809_/B _14809_/Y _14817_/X VGND VGND VPWR VPWR _14818_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15798_ _15670_/X _15797_/Y _15670_/X _15797_/Y VGND VGND VPWR VPWR _16217_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14749_ _14749_/A VGND VGND VPWR VPWR _15181_/A sky130_fd_sc_hd__buf_1
XFILLER_32_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08270_ input11/X VGND VGND VPWR VPWR _08363_/B sky130_fd_sc_hd__inv_2
X_16419_ _16474_/Q _16419_/B VGND VGND VPWR VPWR _16429_/B sky130_fd_sc_hd__or2_1
XFILLER_106_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09724_ _09970_/A _09722_/Y _09723_/Y VGND VGND VPWR VPWR _09770_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09655_ _09609_/Y _09653_/X _09654_/Y VGND VGND VPWR VPWR _09655_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08606_ _08605_/X _08417_/Y _08605_/X _08417_/Y VGND VGND VPWR VPWR _08609_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09586_ _09488_/A _09488_/B _09488_/Y VGND VGND VPWR VPWR _09586_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08537_ _08692_/A _10119_/B VGND VGND VPWR VPWR _08876_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08468_ _08505_/B _08464_/Y _08704_/B VGND VGND VPWR VPWR _08468_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10430_ _11791_/A _10430_/B VGND VGND VPWR VPWR _10430_/X sky130_fd_sc_hd__and2_1
X_08399_ _08399_/A _08399_/B VGND VGND VPWR VPWR _08662_/B sky130_fd_sc_hd__or2_1
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10361_ _09975_/A _09975_/B _09975_/Y VGND VGND VPWR VPWR _10362_/A sky130_fd_sc_hd__o21ai_1
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13080_ _13080_/A _13018_/X VGND VGND VPWR VPWR _13080_/X sky130_fd_sc_hd__or2b_1
X_12100_ _12161_/A _12099_/Y _12161_/A _12099_/Y VGND VGND VPWR VPWR _12158_/B sky130_fd_sc_hd__a2bb2o_1
X_10292_ _10213_/A _10213_/B _10213_/Y VGND VGND VPWR VPWR _12704_/A sky130_fd_sc_hd__o21ai_2
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12031_ _12053_/A VGND VGND VPWR VPWR _13188_/A sky130_fd_sc_hd__buf_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13982_ _13863_/X _13981_/Y _13879_/Y VGND VGND VPWR VPWR _13982_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15721_ _15728_/A _15721_/B VGND VGND VPWR VPWR _16119_/A sky130_fd_sc_hd__or2_1
XFILLER_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12933_ _12895_/Y _12931_/X _12932_/Y VGND VGND VPWR VPWR _12933_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15652_ _15651_/A _15650_/Y _15651_/Y _15650_/A _15571_/A VGND VGND VPWR VPWR _16030_/A
+ sky130_fd_sc_hd__a221o_1
X_12864_ _15171_/A _12863_/B _12863_/Y VGND VGND VPWR VPWR _12864_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15583_ _15583_/A _14396_/X VGND VGND VPWR VPWR _15583_/X sky130_fd_sc_hd__or2b_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _15187_/A _14604_/B VGND VGND VPWR VPWR _14605_/A sky130_fd_sc_hd__and2_1
X_12795_ _12858_/A _12858_/B VGND VGND VPWR VPWR _12795_/Y sky130_fd_sc_hd__nor2_1
X_11815_ _11847_/B _11814_/Y _11847_/B _11814_/Y VGND VGND VPWR VPWR _11845_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _14525_/X _14533_/X _14525_/X _14533_/X VGND VGND VPWR VPWR _14536_/B sky130_fd_sc_hd__a2bb2o_1
X_11746_ _11745_/A _11745_/B _10224_/B _11745_/X VGND VGND VPWR VPWR _11747_/A sky130_fd_sc_hd__a22o_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16204_ _16098_/X _16203_/X _16098_/X _16203_/X VGND VGND VPWR VPWR _16205_/B sky130_fd_sc_hd__o2bb2a_1
X_11677_ _11674_/Y _11676_/X _11674_/Y _11676_/X VGND VGND VPWR VPWR _11677_/X sky130_fd_sc_hd__a2bb2o_2
X_14465_ _14465_/A _14465_/B VGND VGND VPWR VPWR _14465_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14396_ _15966_/A _14396_/B VGND VGND VPWR VPWR _14396_/X sky130_fd_sc_hd__or2_1
X_13416_ _14908_/A _13416_/B VGND VGND VPWR VPWR _14351_/B sky130_fd_sc_hd__or2_1
X_10628_ _10628_/A VGND VGND VPWR VPWR _11892_/A sky130_fd_sc_hd__buf_1
XFILLER_127_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16135_ _16388_/A _16135_/B VGND VGND VPWR VPWR _16136_/B sky130_fd_sc_hd__or2_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13347_ _13274_/A _13274_/B _13274_/Y VGND VGND VPWR VPWR _13347_/Y sky130_fd_sc_hd__o21ai_1
X_10559_ _10559_/A VGND VGND VPWR VPWR _11920_/A sky130_fd_sc_hd__inv_2
X_16066_ _16045_/X _16065_/Y _16045_/X _16065_/Y VGND VGND VPWR VPWR _16114_/B sky130_fd_sc_hd__a2bb2o_1
X_13278_ _13278_/A VGND VGND VPWR VPWR _13278_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12229_ _12136_/X _12228_/X _12136_/X _12228_/X VGND VGND VPWR VPWR _12230_/B sky130_fd_sc_hd__a2bb2o_1
X_15017_ _11811_/X _15001_/X _11811_/X _15001_/X VGND VGND VPWR VPWR _15036_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15919_ _15902_/A _15902_/B _15902_/Y VGND VGND VPWR VPWR _15919_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09440_ _09430_/A _09430_/B _09430_/X _09439_/X VGND VGND VPWR VPWR _09440_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09371_ _09430_/B _09371_/B VGND VGND VPWR VPWR _09371_/X sky130_fd_sc_hd__or2_1
X_08322_ _08322_/A _08322_/B VGND VGND VPWR VPWR _08323_/A sky130_fd_sc_hd__or2_1
XFILLER_60_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08253_ input33/X VGND VGND VPWR VPWR _08254_/B sky130_fd_sc_hd__inv_2
XFILLER_20_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09707_ _09707_/A _09707_/B VGND VGND VPWR VPWR _09707_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09638_ _09539_/A _09539_/B _09539_/X VGND VGND VPWR VPWR _09638_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_82_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09569_ _09569_/A _09569_/B VGND VGND VPWR VPWR _09569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12580_ _12580_/A VGND VGND VPWR VPWR _12580_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11600_ _11599_/A _11599_/B _11599_/Y _10982_/X VGND VGND VPWR VPWR _11616_/A sky130_fd_sc_hd__o211a_1
X_11531_ _11519_/X _11530_/Y _11519_/X _11530_/Y VGND VGND VPWR VPWR _11620_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14250_ _14372_/A _15885_/A VGND VGND VPWR VPWR _14250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11462_ _11569_/A _11462_/B VGND VGND VPWR VPWR _12407_/A sky130_fd_sc_hd__or2_1
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14181_ _13442_/A _14127_/A _14125_/Y VGND VGND VPWR VPWR _14181_/Y sky130_fd_sc_hd__a21oi_1
X_13201_ _13153_/Y _13199_/X _13200_/Y VGND VGND VPWR VPWR _13201_/X sky130_fd_sc_hd__o21a_1
X_10413_ _11783_/A _10338_/B _11783_/A _10338_/B VGND VGND VPWR VPWR _10413_/X sky130_fd_sc_hd__a2bb2o_1
X_11393_ _11393_/A VGND VGND VPWR VPWR _11393_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13132_ _15433_/A VGND VGND VPWR VPWR _14068_/A sky130_fd_sc_hd__inv_2
X_10344_ _12605_/A _10344_/B VGND VGND VPWR VPWR _10421_/A sky130_fd_sc_hd__or2_1
XFILLER_124_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13063_ _13063_/A VGND VGND VPWR VPWR _13769_/A sky130_fd_sc_hd__inv_2
X_10275_ _11724_/A VGND VGND VPWR VPWR _12706_/A sky130_fd_sc_hd__buf_1
XFILLER_3_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ _13198_/A _12063_/B VGND VGND VPWR VPWR _12014_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13965_ _13495_/A _13495_/B _13495_/X VGND VGND VPWR VPWR _13965_/X sky130_fd_sc_hd__o21ba_1
XFILLER_19_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15704_ _15991_/A _15825_/B _15703_/Y VGND VGND VPWR VPWR _15704_/Y sky130_fd_sc_hd__o21ai_1
X_13896_ _13857_/X _13895_/Y _13857_/X _13895_/Y VGND VGND VPWR VPWR _13958_/B sky130_fd_sc_hd__a2bb2o_1
X_12916_ _12916_/A VGND VGND VPWR VPWR _12916_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15635_ _16034_/A VGND VGND VPWR VPWR _15671_/A sky130_fd_sc_hd__inv_2
XFILLER_64_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12847_ _12813_/Y _12845_/X _12846_/Y VGND VGND VPWR VPWR _12847_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _15289_/A _15289_/B _15289_/Y _15354_/X VGND VGND VPWR VPWR _15566_/X sky130_fd_sc_hd__o2bb2a_1
X_12778_ _12738_/Y _12776_/X _12777_/Y VGND VGND VPWR VPWR _12778_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15497_ _15548_/A _15548_/B VGND VGND VPWR VPWR _15497_/X sky130_fd_sc_hd__and2_1
X_14517_ _14553_/A _14515_/X _14516_/X VGND VGND VPWR VPWR _14517_/X sky130_fd_sc_hd__o21a_1
X_11729_ _11729_/A VGND VGND VPWR VPWR _11731_/A sky130_fd_sc_hd__inv_2
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14448_ _14465_/A _14465_/B VGND VGND VPWR VPWR _14448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14379_ _14361_/Y _14377_/X _14378_/Y VGND VGND VPWR VPWR _14379_/X sky130_fd_sc_hd__o21a_1
X_16118_ _16050_/X _16117_/Y _16050_/X _16117_/Y VGND VGND VPWR VPWR _16147_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16049_ _15966_/A _15966_/B _15966_/Y VGND VGND VPWR VPWR _16049_/Y sky130_fd_sc_hd__o21ai_1
X_08940_ _08679_/A _08679_/B _08679_/A _08679_/B VGND VGND VPWR VPWR _08940_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08871_ _08871_/A _08871_/B VGND VGND VPWR VPWR _08871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09423_ _09769_/A _09424_/B VGND VGND VPWR VPWR _09423_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09354_ _09354_/A VGND VGND VPWR VPWR _09354_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08305_ _08239_/Y _08296_/A _08239_/A _08296_/Y _08304_/X VGND VGND VPWR VPWR _08505_/B
+ sky130_fd_sc_hd__o221a_1
X_09285_ _09239_/X _09284_/X _09239_/X _09284_/X VGND VGND VPWR VPWR _09286_/A sky130_fd_sc_hd__a2bb2o_1
X_08236_ input7/X VGND VGND VPWR VPWR _08237_/A sky130_fd_sc_hd__inv_2
XFILLER_119_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10060_ _10059_/A _10059_/B _10216_/A _10059_/Y VGND VGND VPWR VPWR _10063_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_125_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13750_ _13757_/A _13757_/B VGND VGND VPWR VPWR _13750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10962_ _10962_/A _11997_/A VGND VGND VPWR VPWR _10962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12701_ _12701_/A VGND VGND VPWR VPWR _12703_/A sky130_fd_sc_hd__buf_1
X_15420_ _15420_/A _15420_/B VGND VGND VPWR VPWR _15420_/X sky130_fd_sc_hd__or2_1
X_13681_ _14505_/A VGND VGND VPWR VPWR _13684_/A sky130_fd_sc_hd__inv_2
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10893_ _10893_/A VGND VGND VPWR VPWR _10893_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12632_ _14190_/A _12630_/X _12631_/X VGND VGND VPWR VPWR _12632_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12563_ _12625_/A _12625_/B VGND VGND VPWR VPWR _14208_/A sky130_fd_sc_hd__and2_1
X_15351_ _15351_/A _15351_/B VGND VGND VPWR VPWR _15351_/X sky130_fd_sc_hd__or2_1
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14302_ _13443_/X _14301_/X _13443_/X _14301_/X VGND VGND VPWR VPWR _14303_/B sky130_fd_sc_hd__a2bb2oi_1
X_12494_ _12494_/A _12494_/B VGND VGND VPWR VPWR _12494_/Y sky130_fd_sc_hd__nand2_1
X_15282_ _14746_/A _15240_/B _15240_/Y _15281_/X VGND VGND VPWR VPWR _15282_/X sky130_fd_sc_hd__a2bb2o_1
X_11514_ _12373_/A VGND VGND VPWR VPWR _12684_/A sky130_fd_sc_hd__buf_1
X_14233_ _12616_/A _14232_/X _12616_/A _14232_/X VGND VGND VPWR VPWR _14251_/B sky130_fd_sc_hd__a2bb2o_1
X_11445_ _12344_/A VGND VGND VPWR VPWR _15534_/A sky130_fd_sc_hd__buf_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14164_ _12641_/A _14163_/X _12641_/A _14163_/X VGND VGND VPWR VPWR _14166_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11376_ _11258_/X _11375_/Y _11258_/X _11375_/Y VGND VGND VPWR VPWR _11377_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14095_ _14051_/X _14094_/X _14051_/X _14094_/X VGND VGND VPWR VPWR _14095_/Y sky130_fd_sc_hd__a2bb2oi_1
X_13115_ _15249_/A _13115_/B VGND VGND VPWR VPWR _13115_/Y sky130_fd_sc_hd__nand2_1
X_10327_ _10295_/X _10326_/X _10295_/X _10326_/X VGND VGND VPWR VPWR _10328_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13031_/X _13045_/X _13031_/X _13045_/X VGND VGND VPWR VPWR _13123_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _09269_/B _10243_/B _10243_/X _10688_/A VGND VGND VPWR VPWR _10826_/A sky130_fd_sc_hd__a22o_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10189_ _10241_/B _10151_/B _10151_/Y _10973_/A VGND VGND VPWR VPWR _11148_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_94_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14997_ _11713_/A _11720_/B _10521_/A _11713_/Y VGND VGND VPWR VPWR _14997_/X sky130_fd_sc_hd__o2bb2a_1
X_13948_ _15406_/A _13948_/B VGND VGND VPWR VPWR _13948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13879_ _13879_/A _13981_/B VGND VGND VPWR VPWR _13879_/Y sky130_fd_sc_hd__nand2_1
X_15618_ _15616_/A _15617_/A _15616_/Y _15617_/Y _15595_/A VGND VGND VPWR VPWR _16038_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15549_ _15497_/X _15547_/X _15579_/B VGND VGND VPWR VPWR _15549_/X sky130_fd_sc_hd__o21a_1
X_09070_ _09070_/A _09070_/B VGND VGND VPWR VPWR _09071_/B sky130_fd_sc_hd__or2_1
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09972_ _09972_/A _09972_/B VGND VGND VPWR VPWR _09972_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08923_ _09293_/B VGND VGND VPWR VPWR _10228_/B sky130_fd_sc_hd__inv_2
XFILLER_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08854_ _08937_/B VGND VGND VPWR VPWR _09041_/B sky130_fd_sc_hd__inv_2
XFILLER_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08785_ _10012_/A VGND VGND VPWR VPWR _09470_/A sky130_fd_sc_hd__buf_1
XFILLER_80_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09406_ _09407_/A _09407_/B VGND VGND VPWR VPWR _10892_/A sky130_fd_sc_hd__and2_1
X_09337_ _08770_/A _08768_/Y _10038_/A _09336_/X VGND VGND VPWR VPWR _09337_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09268_ _10243_/A VGND VGND VPWR VPWR _09269_/B sky130_fd_sc_hd__buf_1
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09199_ _09199_/A VGND VGND VPWR VPWR _09199_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11230_ _12224_/A _11230_/B VGND VGND VPWR VPWR _11230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11161_ _11131_/X _11160_/X _11131_/X _11160_/X VGND VGND VPWR VPWR _11302_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10112_ _10112_/A _10112_/B VGND VGND VPWR VPWR _10113_/A sky130_fd_sc_hd__or2_1
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11092_ _11195_/A _11090_/X _11091_/X VGND VGND VPWR VPWR _11092_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14920_ _15544_/A _14920_/B VGND VGND VPWR VPWR _14920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10043_ _10043_/A _10083_/B VGND VGND VPWR VPWR _10043_/X sky130_fd_sc_hd__and2_1
X_14851_ _14953_/A _14953_/B VGND VGND VPWR VPWR _14851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13802_ _13774_/X _13801_/X _13774_/X _13801_/X VGND VGND VPWR VPWR _13858_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14782_ _14782_/A _14782_/B VGND VGND VPWR VPWR _14782_/X sky130_fd_sc_hd__and2_1
XFILLER_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11994_ _11994_/A VGND VGND VPWR VPWR _12082_/B sky130_fd_sc_hd__inv_2
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13733_ _13733_/A _13697_/X VGND VGND VPWR VPWR _13733_/X sky130_fd_sc_hd__or2b_1
X_10945_ _10944_/Y _10790_/X _10836_/Y VGND VGND VPWR VPWR _10945_/X sky130_fd_sc_hd__o21a_1
X_16452_ _16432_/X _16444_/Y _16450_/X _16451_/X VGND VGND VPWR VPWR _16472_/D sky130_fd_sc_hd__o211ai_4
X_13664_ _13697_/A _13697_/B VGND VGND VPWR VPWR _13733_/A sky130_fd_sc_hd__and2_1
X_10876_ _10876_/A _09412_/X VGND VGND VPWR VPWR _10877_/A sky130_fd_sc_hd__or2b_1
X_16383_ _08230_/A _16458_/Q _08233_/A _16396_/C _16343_/A VGND VGND VPWR VPWR _16458_/D
+ sky130_fd_sc_hd__o221a_2
X_12615_ _14235_/A _14235_/B VGND VGND VPWR VPWR _12616_/A sky130_fd_sc_hd__nand2_1
X_15403_ _15462_/A _15401_/X _15402_/X VGND VGND VPWR VPWR _15403_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15334_ _15387_/A _15332_/X _15333_/X VGND VGND VPWR VPWR _15334_/X sky130_fd_sc_hd__o21a_1
X_13595_ _13578_/X _13594_/Y _13578_/X _13594_/Y VGND VGND VPWR VPWR _13630_/B sky130_fd_sc_hd__a2bb2o_1
X_12546_ _14916_/A _11453_/B _11453_/Y VGND VGND VPWR VPWR _12547_/A sky130_fd_sc_hd__o21ai_1
X_12477_ _12402_/A _12357_/X _12401_/X VGND VGND VPWR VPWR _12477_/Y sky130_fd_sc_hd__o21ai_1
X_15265_ _15211_/A _15211_/B _15211_/Y VGND VGND VPWR VPWR _15265_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14216_ _15872_/A _14260_/B VGND VGND VPWR VPWR _14216_/Y sky130_fd_sc_hd__nor2_1
X_11428_ _11252_/X _11427_/Y _11252_/X _11427_/Y VGND VGND VPWR VPWR _12585_/A sky130_fd_sc_hd__a2bb2o_1
X_15196_ _15196_/A _15196_/B VGND VGND VPWR VPWR _15196_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_4 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11359_ _11569_/A _11359_/B VGND VGND VPWR VPWR _12303_/A sky130_fd_sc_hd__or2_1
X_14147_ _14147_/A _14068_/X VGND VGND VPWR VPWR _14147_/X sky130_fd_sc_hd__or2b_1
XFILLER_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14078_ _14055_/X _14077_/X _14055_/X _14077_/X VGND VGND VPWR VPWR _14115_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _13055_/A _13027_/X _13028_/X VGND VGND VPWR VPWR _13029_/X sky130_fd_sc_hd__o21a_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer27 _16231_/B VGND VGND VPWR VPWR _16318_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08570_ _08713_/B VGND VGND VPWR VPWR _08572_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer16 rebuffer17/X VGND VGND VPWR VPWR rebuffer16/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09122_ _09122_/A VGND VGND VPWR VPWR _09122_/Y sky130_fd_sc_hd__inv_2
X_09053_ _08711_/Y _09052_/Y _08737_/X VGND VGND VPWR VPWR _09054_/A sky130_fd_sc_hd__o21ai_1
XFILLER_104_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09955_ _09955_/A _09955_/B VGND VGND VPWR VPWR _09955_/X sky130_fd_sc_hd__and2_1
XFILLER_131_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09886_/A _09886_/B VGND VGND VPWR VPWR _09887_/B sky130_fd_sc_hd__or2_1
X_08906_ _08905_/Y _08861_/X _08905_/Y _08861_/X VGND VGND VPWR VPWR _08972_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _09459_/A VGND VGND VPWR VPWR _09502_/A sky130_fd_sc_hd__buf_1
XFILLER_18_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08768_ _08770_/B VGND VGND VPWR VPWR _08768_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08699_ _08699_/A VGND VGND VPWR VPWR _08699_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10730_ _09960_/A _09645_/B _09645_/Y VGND VGND VPWR VPWR _10732_/A sky130_fd_sc_hd__o21ai_1
XFILLER_40_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10661_ _10660_/A _10660_/B _10660_/Y _09393_/A VGND VGND VPWR VPWR _10795_/A sky130_fd_sc_hd__o211a_1
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12400_ _13545_/A _12401_/B VGND VGND VPWR VPWR _12402_/A sky130_fd_sc_hd__and2_1
XFILLER_9_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13380_ _13370_/X _13379_/X _13370_/X _13379_/X VGND VGND VPWR VPWR _13446_/B sky130_fd_sc_hd__a2bb2o_1
X_10592_ _11841_/A _10531_/B _10531_/Y VGND VGND VPWR VPWR _10592_/Y sky130_fd_sc_hd__o21ai_1
X_12331_ _12575_/A _12334_/B VGND VGND VPWR VPWR _12331_/Y sky130_fd_sc_hd__nor2_1
X_12262_ _12262_/A VGND VGND VPWR VPWR _12262_/Y sky130_fd_sc_hd__inv_2
X_15050_ _15051_/A _15051_/B VGND VGND VPWR VPWR _15052_/A sky130_fd_sc_hd__and2_1
XFILLER_5_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11213_ _11213_/A _11219_/B VGND VGND VPWR VPWR _13334_/A sky130_fd_sc_hd__or2_1
X_14001_ _13995_/A _13995_/B _13995_/Y VGND VGND VPWR VPWR _14001_/Y sky130_fd_sc_hd__o21ai_1
X_12193_ _12252_/A _12252_/B VGND VGND VPWR VPWR _12193_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11144_ _11604_/A _11144_/B VGND VGND VPWR VPWR _11145_/A sky130_fd_sc_hd__or2_1
XFILLER_1_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15952_ _15952_/A _15952_/B VGND VGND VPWR VPWR _15952_/X sky130_fd_sc_hd__or2_1
X_11075_ _12137_/A VGND VGND VPWR VPWR _15392_/A sky130_fd_sc_hd__buf_1
XFILLER_49_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14903_ _14047_/X _14902_/X _14047_/X _14902_/X VGND VGND VPWR VPWR _14904_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10026_ _09324_/A _08793_/B _10047_/B _10025_/X VGND VGND VPWR VPWR _10026_/X sky130_fd_sc_hd__o22a_1
X_15883_ _15886_/A _15886_/B VGND VGND VPWR VPWR _15883_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14834_ _14747_/X _14833_/Y _14764_/Y VGND VGND VPWR VPWR _14834_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14765_ _14833_/A _14833_/B _14764_/Y VGND VGND VPWR VPWR _14765_/Y sky130_fd_sc_hd__o21ai_1
X_11977_ _11939_/Y _11975_/X _11976_/Y VGND VGND VPWR VPWR _11977_/X sky130_fd_sc_hd__o21a_1
X_10928_ _12104_/A VGND VGND VPWR VPWR _11002_/A sky130_fd_sc_hd__inv_2
X_13716_ _13716_/A _13779_/B VGND VGND VPWR VPWR _13716_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16435_ _16462_/Q _16461_/Q _16464_/Q _16463_/Q VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__or4_1
X_14696_ _14737_/A _14737_/B VGND VGND VPWR VPWR _14784_/A sky130_fd_sc_hd__and2_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10859_ _10915_/A _10916_/B VGND VGND VPWR VPWR _11025_/A sky130_fd_sc_hd__and2_1
X_13647_ _15044_/A _13507_/B _13507_/Y VGND VGND VPWR VPWR _13647_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16366_ _16326_/A _16326_/B _16326_/Y VGND VGND VPWR VPWR _16366_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _12844_/A _13560_/B _13561_/Y _13577_/X VGND VGND VPWR VPWR _13578_/X sky130_fd_sc_hd__o22a_1
X_16297_ _16260_/A _16326_/A _16260_/Y VGND VGND VPWR VPWR _16297_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_117_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12529_ _13440_/A _11377_/B _11377_/Y VGND VGND VPWR VPWR _12530_/B sky130_fd_sc_hd__o21a_1
X_15317_ _15337_/A _15337_/B VGND VGND VPWR VPWR _15381_/A sky130_fd_sc_hd__and2_1
XFILLER_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15248_ _15223_/X _15247_/Y _15223_/X _15247_/Y VGND VGND VPWR VPWR _15249_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15179_ _15113_/A _15113_/B _15113_/Y VGND VGND VPWR VPWR _15179_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09740_ _09740_/A _09740_/B VGND VGND VPWR VPWR _09743_/B sky130_fd_sc_hd__or2_1
.ends

