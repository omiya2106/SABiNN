* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt user_project_wrapper VGND VPWR wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09671_ _10763_/A VGND VGND VPWR VPWR _09672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08622_ _08622_/A VGND VGND VPWR VPWR _10112_/B sky130_fd_sc_hd__inv_2
XFILLER_54_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08553_ _09470_/B VGND VGND VPWR VPWR _08688_/A sky130_fd_sc_hd__buf_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08484_ _08275_/A _08357_/B _08480_/Y _08483_/X VGND VGND VPWR VPWR _08625_/A sky130_fd_sc_hd__o22a_1
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09105_ _08674_/Y _09028_/A _09030_/B VGND VGND VPWR VPWR _09105_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09036_ _09555_/B _09036_/B VGND VGND VPWR VPWR _09037_/B sky130_fd_sc_hd__or2_1
XFILLER_117_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09938_ _09936_/X _09937_/Y _09791_/C _09874_/X _09888_/X VGND VGND VPWR VPWR _09938_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09869_ _09451_/Y _09868_/X _09472_/X VGND VGND VPWR VPWR _09869_/X sky130_fd_sc_hd__o21a_1
XFILLER_73_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11900_ _11900_/A VGND VGND VPWR VPWR _11900_/Y sky130_fd_sc_hd__inv_2
X_12880_ _14599_/A _12942_/B VGND VGND VPWR VPWR _12880_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11831_ _11790_/A _11790_/B _11790_/Y VGND VGND VPWR VPWR _11831_/X sky130_fd_sc_hd__a21o_1
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14581_/A _14581_/B VGND VGND VPWR VPWR _14550_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13503_/A VGND VGND VPWR VPWR _15046_/A sky130_fd_sc_hd__buf_1
X_11762_ _11762_/A _11762_/B VGND VGND VPWR VPWR _11762_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14468_/A _14468_/B _14468_/Y VGND VGND VPWR VPWR _14481_/Y sky130_fd_sc_hd__o21ai_1
X_10713_ _11910_/A VGND VGND VPWR VPWR _13696_/A sky130_fd_sc_hd__buf_1
XFILLER_41_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11693_ _12426_/B VGND VGND VPWR VPWR _11694_/B sky130_fd_sc_hd__inv_2
X_16220_ _16253_/B VGND VGND VPWR VPWR _16320_/A sky130_fd_sc_hd__clkbuf_2
X_13432_ _14111_/A _13435_/B VGND VGND VPWR VPWR _13432_/Y sky130_fd_sc_hd__nor2_1
X_10644_ _10644_/A VGND VGND VPWR VPWR _10644_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16151_ _15818_/X _16150_/X _15818_/X _16150_/X VGND VGND VPWR VPWR _16152_/B sky130_fd_sc_hd__a2bb2o_1
X_13363_ _13390_/A _13361_/X _13362_/X VGND VGND VPWR VPWR _13363_/X sky130_fd_sc_hd__o21a_1
X_10575_ _10675_/A _12695_/A _10574_/Y VGND VGND VPWR VPWR _10575_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12314_ _12314_/A _12314_/B VGND VGND VPWR VPWR _12314_/Y sky130_fd_sc_hd__nand2_1
X_15102_ _12383_/Y _15101_/X _12383_/Y _15101_/X VGND VGND VPWR VPWR _15104_/B sky130_fd_sc_hd__a2bb2o_1
Xrebuffer7 rebuffer8/X VGND VGND VPWR VPWR rebuffer7/X sky130_fd_sc_hd__dlygate4sd1_1
X_16082_ _16084_/A _16084_/B VGND VGND VPWR VPWR _16082_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13294_ _14736_/A _13294_/B VGND VGND VPWR VPWR _13294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12245_ _14023_/A _12217_/B _12217_/Y _12244_/X VGND VGND VPWR VPWR _12245_/X sky130_fd_sc_hd__a2bb2o_1
X_15033_ _15076_/A _15031_/X _15032_/X VGND VGND VPWR VPWR _15033_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12176_ _12176_/A _12176_/B VGND VGND VPWR VPWR _12176_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11127_ _12189_/A VGND VGND VPWR VPWR _13715_/A sky130_fd_sc_hd__buf_1
X_15935_ _15891_/X _15934_/Y _15891_/X _15934_/Y VGND VGND VPWR VPWR _15954_/B sky130_fd_sc_hd__a2bb2o_1
X_11058_ _10911_/X _11057_/Y _10911_/X _11057_/Y VGND VGND VPWR VPWR _11078_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15866_ _15866_/A VGND VGND VPWR VPWR _15896_/A sky130_fd_sc_hd__inv_2
XFILLER_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10009_ _10009_/A _10009_/B VGND VGND VPWR VPWR _10035_/B sky130_fd_sc_hd__nor2_1
X_14817_ _14812_/A _14812_/B _14812_/Y _14816_/X VGND VGND VPWR VPWR _14817_/X sky130_fd_sc_hd__o2bb2a_1
X_15797_ _16099_/A _15800_/B VGND VGND VPWR VPWR _15797_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14748_ _14667_/X _14681_/A _14680_/X VGND VGND VPWR VPWR _14748_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14679_ _15184_/A _14680_/B VGND VGND VPWR VPWR _14681_/A sky130_fd_sc_hd__and2_1
XFILLER_60_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16418_ _16473_/Q VGND VGND VPWR VPWR _16419_/B sky130_fd_sc_hd__inv_2
XFILLER_32_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16349_ _16335_/X _16348_/Y _16335_/X _16348_/Y VGND VGND VPWR VPWR _16349_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09723_ _09723_/A _09723_/B VGND VGND VPWR VPWR _09723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09654_ _09981_/A _09654_/B VGND VGND VPWR VPWR _09654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08605_ _09249_/A _09217_/B _10015_/A _08604_/Y VGND VGND VPWR VPWR _08605_/X sky130_fd_sc_hd__o22a_1
XFILLER_70_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09585_ _09993_/A _09662_/B VGND VGND VPWR VPWR _09585_/Y sky130_fd_sc_hd__nor2_1
X_08536_ _08535_/A _08453_/Y _08535_/Y _08453_/A VGND VGND VPWR VPWR _10119_/B sky130_fd_sc_hd__o22a_1
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08467_ _09146_/A VGND VGND VPWR VPWR _08704_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08398_ _08398_/A VGND VGND VPWR VPWR _08398_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10360_ _13524_/A _10319_/B _10319_/X _10359_/X VGND VGND VPWR VPWR _10360_/X sky130_fd_sc_hd__o22a_1
X_10291_ _12707_/A _10291_/B VGND VGND VPWR VPWR _10291_/X sky130_fd_sc_hd__or2_1
X_09019_ _09019_/A VGND VGND VPWR VPWR _09531_/B sky130_fd_sc_hd__inv_2
X_12030_ _13078_/A _11972_/B _11972_/Y VGND VGND VPWR VPWR _12030_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13981_ _13862_/X _13980_/Y _13878_/Y VGND VGND VPWR VPWR _13981_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15720_ _14923_/X _15719_/X _14923_/X _15719_/X VGND VGND VPWR VPWR _15721_/B sky130_fd_sc_hd__a2bb2oi_1
X_12932_ _12932_/A _12932_/B VGND VGND VPWR VPWR _12932_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15651_ _15651_/A VGND VGND VPWR VPWR _15651_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14602_ _15187_/A _14603_/B VGND VGND VPWR VPWR _14604_/A sky130_fd_sc_hd__and2_1
XFILLER_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12863_ _12790_/X _12862_/X _12790_/X _12862_/X VGND VGND VPWR VPWR _12864_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15582_ _16051_/A VGND VGND VPWR VPWR _15685_/A sky130_fd_sc_hd__inv_2
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12784_/A _12784_/B _12784_/Y VGND VGND VPWR VPWR _12794_/Y sky130_fd_sc_hd__o21ai_1
X_11814_ _11812_/X _11814_/B VGND VGND VPWR VPWR _11814_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14524_/X _14532_/X _14524_/X _14532_/X VGND VGND VPWR VPWR _14535_/B sky130_fd_sc_hd__a2bb2o_1
X_11745_ _11745_/A _11745_/B VGND VGND VPWR VPWR _11745_/X sky130_fd_sc_hd__or2_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ _14464_/A _14464_/B VGND VGND VPWR VPWR _14464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16203_ _16099_/A _16099_/B _16099_/Y VGND VGND VPWR VPWR _16203_/X sky130_fd_sc_hd__o21a_1
X_13415_ _14908_/A _13415_/B VGND VGND VPWR VPWR _14350_/B sky130_fd_sc_hd__or2_1
X_11676_ _15554_/A _11676_/B VGND VGND VPWR VPWR _12643_/B sky130_fd_sc_hd__or2_1
X_14395_ _15966_/A _14395_/B VGND VGND VPWR VPWR _15583_/B sky130_fd_sc_hd__or2_1
X_10627_ _12043_/A VGND VGND VPWR VPWR _15212_/B sky130_fd_sc_hd__inv_2
X_16134_ _16122_/X _16133_/X _16122_/X _16133_/X VGND VGND VPWR VPWR _16135_/B sky130_fd_sc_hd__a2bb2o_1
X_13346_ _13274_/A _13274_/B _13274_/Y VGND VGND VPWR VPWR _13346_/Y sky130_fd_sc_hd__o21ai_1
X_10558_ _09421_/A _09126_/B _09126_/Y VGND VGND VPWR VPWR _10558_/X sky130_fd_sc_hd__o21a_1
X_16065_ _16046_/A _16046_/B _16046_/Y VGND VGND VPWR VPWR _16065_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_115_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13277_ _13264_/Y _13275_/X _13276_/Y VGND VGND VPWR VPWR _13278_/A sky130_fd_sc_hd__o21ai_2
X_12228_ _12140_/X _12227_/X _12140_/X _12227_/X VGND VGND VPWR VPWR _12229_/B sky130_fd_sc_hd__a2bb2o_1
X_15016_ _15038_/A _15038_/B VGND VGND VPWR VPWR _15067_/A sky130_fd_sc_hd__and2_1
X_10489_ _10489_/A VGND VGND VPWR VPWR _10489_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12159_ _12198_/A VGND VGND VPWR VPWR _13202_/A sky130_fd_sc_hd__buf_1
XFILLER_96_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15918_ _15970_/A _15970_/B VGND VGND VPWR VPWR _15918_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15849_ _14183_/A _15848_/X _12634_/X VGND VGND VPWR VPWR _15849_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09370_ _09430_/B _09370_/B VGND VGND VPWR VPWR _09370_/X sky130_fd_sc_hd__or2_1
X_08321_ _08321_/A input19/X VGND VGND VPWR VPWR _08322_/B sky130_fd_sc_hd__nor2_1
X_08252_ input17/X VGND VGND VPWR VPWR _08326_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_20_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09706_ _09689_/A _09689_/B _09692_/A VGND VGND VPWR VPWR _09963_/A sky130_fd_sc_hd__a21bo_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09637_ _09958_/A _09640_/B VGND VGND VPWR VPWR _09637_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09568_ _09560_/X _09567_/X _09560_/X _09567_/X VGND VGND VPWR VPWR _09569_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08519_ _09525_/A VGND VGND VPWR VPWR _09476_/B sky130_fd_sc_hd__inv_2
XFILLER_70_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11530_ _11615_/B VGND VGND VPWR VPWR _11531_/B sky130_fd_sc_hd__inv_2
XFILLER_11_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09499_ _08831_/X _09463_/X _08831_/X _09463_/X VGND VGND VPWR VPWR _09500_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_109_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11461_ _14137_/A _11358_/B _11358_/Y _12508_/A VGND VGND VPWR VPWR _11569_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14180_ _13441_/A _14126_/A _14124_/Y VGND VGND VPWR VPWR _14180_/Y sky130_fd_sc_hd__a21oi_1
X_13200_ _13200_/A _13200_/B VGND VGND VPWR VPWR _13200_/Y sky130_fd_sc_hd__nand2_1
X_10412_ _09296_/Y _10411_/Y _09296_/A _10411_/A _09391_/A VGND VGND VPWR VPWR _12826_/A
+ sky130_fd_sc_hd__o221a_2
X_11392_ _08969_/X _11391_/X _08969_/X _11391_/X VGND VGND VPWR VPWR _11393_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_124_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13131_ _14148_/A VGND VGND VPWR VPWR _13449_/A sky130_fd_sc_hd__buf_1
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10343_ _10352_/A _10342_/X _10352_/A _10342_/X VGND VGND VPWR VPWR _10355_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13062_ _15246_/A _13117_/B VGND VGND VPWR VPWR _13062_/Y sky130_fd_sc_hd__nor2_1
X_10274_ _11732_/A VGND VGND VPWR VPWR _11727_/A sky130_fd_sc_hd__buf_1
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12013_ _13058_/A _12068_/B VGND VGND VPWR VPWR _12013_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15703_ _15991_/A _15825_/B VGND VGND VPWR VPWR _15703_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13964_ _13494_/A _13494_/B _13494_/X VGND VGND VPWR VPWR _13964_/X sky130_fd_sc_hd__o21ba_1
XFILLER_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13895_ _13856_/X _13894_/Y _13856_/X _13894_/Y VGND VGND VPWR VPWR _13957_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12915_ _12915_/A _12915_/B VGND VGND VPWR VPWR _12915_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15634_ _15632_/A _15633_/A _15632_/Y _15633_/Y _15571_/A VGND VGND VPWR VPWR _16034_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12846_ _12817_/Y _12844_/X _12845_/Y VGND VGND VPWR VPWR _12846_/X sky130_fd_sc_hd__o21a_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _12427_/X _15564_/Y _12427_/X _15564_/Y VGND VGND VPWR VPWR _15565_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14552_/A _14514_/X _14515_/X VGND VGND VPWR VPWR _14516_/X sky130_fd_sc_hd__o21a_1
X_12777_ _12742_/Y _12775_/X _12776_/Y VGND VGND VPWR VPWR _12777_/X sky130_fd_sc_hd__o21a_1
X_15496_ _15483_/X _15495_/X _15483_/X _15495_/X VGND VGND VPWR VPWR _15548_/B sky130_fd_sc_hd__a2bb2o_1
X_11728_ _11727_/A _11733_/A _11727_/Y VGND VGND VPWR VPWR _11728_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11659_ _11583_/X _11658_/Y _11583_/X _11658_/Y VGND VGND VPWR VPWR _11661_/B sky130_fd_sc_hd__a2bb2o_1
X_14447_ _14464_/A _14464_/B VGND VGND VPWR VPWR _14447_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14378_ _14360_/Y _14376_/X _14377_/Y VGND VGND VPWR VPWR _14378_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16117_ _16051_/A _16051_/B _16051_/Y VGND VGND VPWR VPWR _16117_/Y sky130_fd_sc_hd__o21ai_1
X_13329_ _14732_/A _13288_/B _13288_/Y VGND VGND VPWR VPWR _13329_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16048_ _16051_/A _16051_/B VGND VGND VPWR VPWR _16048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08870_ _08986_/A _08986_/B VGND VGND VPWR VPWR _08870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09422_ _09271_/A _09420_/Y _09421_/Y VGND VGND VPWR VPWR _09424_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09353_ _09353_/A VGND VGND VPWR VPWR _09353_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08304_ _08304_/A VGND VGND VPWR VPWR _08304_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09284_ _09238_/X _09283_/X _09238_/X _09283_/X VGND VGND VPWR VPWR _09285_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08235_ input7/X _08235_/B VGND VGND VPWR VPWR _08238_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08999_ _11411_/B VGND VGND VPWR VPWR _11393_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10961_ _12080_/A VGND VGND VPWR VPWR _13506_/A sky130_fd_sc_hd__buf_1
XFILLER_16_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13680_ _14504_/A VGND VGND VPWR VPWR _13683_/A sky130_fd_sc_hd__inv_2
X_12700_ _10310_/Y _12659_/Y _10310_/Y _12659_/Y VGND VGND VPWR VPWR _12701_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_16_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12631_ _14195_/A _12629_/X _12630_/X VGND VGND VPWR VPWR _12631_/X sky130_fd_sc_hd__o21a_1
X_10892_ _13088_/A _10749_/B _10749_/Y VGND VGND VPWR VPWR _10892_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12562_ _14914_/A _12346_/B _12346_/Y VGND VGND VPWR VPWR _12563_/A sky130_fd_sc_hd__o21ai_1
X_15350_ _15363_/A _15348_/X _15349_/X VGND VGND VPWR VPWR _15350_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14301_ _13442_/X _14300_/X _13442_/X _14300_/X VGND VGND VPWR VPWR _14302_/B sky130_fd_sc_hd__a2bb2oi_1
X_12493_ _12487_/Y _12492_/Y _12487_/Y _12492_/Y VGND VGND VPWR VPWR _12496_/B sky130_fd_sc_hd__a2bb2o_1
X_15281_ _14664_/A _15243_/B _15243_/Y _15280_/X VGND VGND VPWR VPWR _15281_/X sky130_fd_sc_hd__a2bb2o_1
X_11513_ _11513_/A _11513_/B VGND VGND VPWR VPWR _11513_/Y sky130_fd_sc_hd__nand2_1
X_14232_ _12617_/A _14231_/Y _12617_/A _14231_/Y VGND VGND VPWR VPWR _14250_/B sky130_fd_sc_hd__a2bb2o_1
X_11444_ _11439_/Y _12566_/A _11443_/Y VGND VGND VPWR VPWR _11449_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14163_ _12642_/A _14162_/X _12642_/A _14162_/X VGND VGND VPWR VPWR _14165_/B sky130_fd_sc_hd__a2bb2o_1
X_11375_ _11393_/A _11375_/B VGND VGND VPWR VPWR _12311_/A sky130_fd_sc_hd__or2_1
XFILLER_125_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14094_ _14050_/X _14093_/X _14050_/X _14093_/X VGND VGND VPWR VPWR _14094_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_79_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13114_ _13072_/Y _13112_/X _13113_/Y VGND VGND VPWR VPWR _13114_/X sky130_fd_sc_hd__o21a_1
X_10326_ _10325_/A _10325_/B _10325_/Y VGND VGND VPWR VPWR _10326_/X sky130_fd_sc_hd__a21o_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13045_ _13045_/A _13033_/X VGND VGND VPWR VPWR _13045_/X sky130_fd_sc_hd__or2b_1
X_10257_ _09274_/B _10244_/B _10244_/X _10571_/A VGND VGND VPWR VPWR _10692_/A sky130_fd_sc_hd__a22o_1
XFILLER_3_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10188_ _10242_/B _10155_/B _10155_/Y _10822_/A VGND VGND VPWR VPWR _10975_/A sky130_fd_sc_hd__o2bb2a_1
X_14996_ _14996_/A _15728_/A VGND VGND VPWR VPWR _16125_/A sky130_fd_sc_hd__or2_1
XFILLER_66_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13947_ _15406_/A _13947_/B VGND VGND VPWR VPWR _13947_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15617_ _15617_/A VGND VGND VPWR VPWR _15617_/Y sky130_fd_sc_hd__clkinvlp_2
X_13878_ _13878_/A _13980_/B VGND VGND VPWR VPWR _13878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12829_ _10623_/A _11719_/A _10521_/A _11720_/B VGND VGND VPWR VPWR _12830_/B sky130_fd_sc_hd__o22a_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15548_ _15548_/A _15548_/B VGND VGND VPWR VPWR _15579_/B sky130_fd_sc_hd__or2_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15479_ _15458_/A _15458_/B _15458_/Y _15478_/X VGND VGND VPWR VPWR _15479_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_30_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09971_ _09971_/A VGND VGND VPWR VPWR _09971_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08922_ _08922_/A _08922_/B VGND VGND VPWR VPWR _09292_/B sky130_fd_sc_hd__nand2_2
XFILLER_111_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08853_ _08916_/A _08913_/B VGND VGND VPWR VPWR _08937_/B sky130_fd_sc_hd__or2_1
XFILLER_111_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08784_ _08786_/B VGND VGND VPWR VPWR _08784_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09405_ _09403_/X _09101_/A _08664_/X _09404_/Y VGND VGND VPWR VPWR _09407_/B sky130_fd_sc_hd__o22a_1
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09336_ _08770_/A _08768_/Y _10038_/A _09335_/X VGND VGND VPWR VPWR _09336_/X sky130_fd_sc_hd__o22a_1
X_09267_ _10243_/A VGND VGND VPWR VPWR _09268_/B sky130_fd_sc_hd__buf_1
XFILLER_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09198_ _09198_/A VGND VGND VPWR VPWR _09198_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11160_ _13503_/A _11306_/B _13503_/A _11306_/B VGND VGND VPWR VPWR _11160_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_134_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11091_ _11204_/A _11089_/X _11090_/X VGND VGND VPWR VPWR _11091_/X sky130_fd_sc_hd__o21a_1
X_10111_ _10111_/A _10111_/B VGND VGND VPWR VPWR _10112_/A sky130_fd_sc_hd__or2_1
XFILLER_88_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10042_ _10027_/X _10041_/Y _10027_/X _10041_/Y VGND VGND VPWR VPWR _10083_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14850_ _14835_/X _14849_/X _14835_/X _14849_/X VGND VGND VPWR VPWR _14953_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14781_ _14737_/X _14780_/X _14737_/X _14780_/X VGND VGND VPWR VPWR _14782_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13801_ _13773_/X _13800_/Y _13773_/X _13800_/Y VGND VGND VPWR VPWR _13857_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13732_ _13732_/A _13696_/X VGND VGND VPWR VPWR _13732_/X sky130_fd_sc_hd__or2b_1
XFILLER_56_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11993_ _11992_/A _11992_/B _11992_/X _11928_/B VGND VGND VPWR VPWR _12082_/B sky130_fd_sc_hd__a22o_1
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10944_ _09967_/Y _10942_/A _10081_/A _10942_/Y _11593_/A VGND VGND VPWR VPWR _12162_/A
+ sky130_fd_sc_hd__a221o_2
X_16451_ _16437_/D _16419_/B _16445_/X _16448_/X VGND VGND VPWR VPWR _16451_/X sky130_fd_sc_hd__o211a_1
X_10875_ _10878_/A VGND VGND VPWR VPWR _14626_/A sky130_fd_sc_hd__buf_1
XFILLER_71_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13663_ _13696_/A _13696_/B VGND VGND VPWR VPWR _13732_/A sky130_fd_sc_hd__and2_1
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16382_ _16312_/Y _16381_/Y _16312_/Y _16381_/Y VGND VGND VPWR VPWR _16396_/C sky130_fd_sc_hd__a2bb2o_1
X_12614_ _12614_/A VGND VGND VPWR VPWR _12614_/Y sky130_fd_sc_hd__clkinvlp_2
X_15402_ _15402_/A _15402_/B VGND VGND VPWR VPWR _15402_/X sky130_fd_sc_hd__or2_1
X_13594_ _13577_/X _13593_/Y _13577_/X _13593_/Y VGND VGND VPWR VPWR _13629_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12545_ _12630_/A _12630_/B VGND VGND VPWR VPWR _14195_/A sky130_fd_sc_hd__and2_1
X_15333_ _15333_/A _15333_/B VGND VGND VPWR VPWR _15333_/X sky130_fd_sc_hd__or2_1
XFILLER_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15264_ _15264_/A _15264_/B VGND VGND VPWR VPWR _15264_/Y sky130_fd_sc_hd__nand2_1
X_12476_ _12466_/X _12476_/B VGND VGND VPWR VPWR _12476_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_125_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14215_ _15872_/A _14259_/B VGND VGND VPWR VPWR _14215_/Y sky130_fd_sc_hd__nor2_1
X_11427_ _14083_/A _11424_/B _11424_/Y _12595_/A VGND VGND VPWR VPWR _11431_/B sky130_fd_sc_hd__o2bb2a_1
X_15195_ _15152_/X _15194_/Y _15152_/X _15194_/Y VGND VGND VPWR VPWR _15196_/B sky130_fd_sc_hd__a2bb2o_1
XANTENNA_5 input33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11358_ _12302_/A _11358_/B VGND VGND VPWR VPWR _11358_/Y sky130_fd_sc_hd__nand2_1
X_14146_ _14002_/X _14146_/B VGND VGND VPWR VPWR _14146_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10309_ _10309_/A _10309_/B VGND VGND VPWR VPWR _10309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14077_ _14054_/X _14076_/X _14054_/X _14076_/X VGND VGND VPWR VPWR _14114_/A sky130_fd_sc_hd__a2bb2o_1
X_11289_ _13043_/A VGND VGND VPWR VPWR _12289_/A sky130_fd_sc_hd__buf_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13028_ _13060_/A _13026_/X _13027_/X VGND VGND VPWR VPWR _13028_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer17 rebuffer18/X VGND VGND VPWR VPWR rebuffer17/X sky130_fd_sc_hd__dlygate4sd1_1
X_14979_ _14977_/Y _14978_/X _14977_/Y _14978_/X VGND VGND VPWR VPWR _14979_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer39 _08372_/X VGND VGND VPWR VPWR _08434_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer28 _08395_/A VGND VGND VPWR VPWR _08934_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09121_ _09549_/B _09033_/B _09034_/B VGND VGND VPWR VPWR _09122_/A sky130_fd_sc_hd__a21bo_1
XFILLER_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09052_ _09052_/A VGND VGND VPWR VPWR _09052_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09954_ _09954_/A VGND VGND VPWR VPWR _09954_/Y sky130_fd_sc_hd__inv_4
XFILLER_58_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _09885_/A _09885_/B VGND VGND VPWR VPWR _09886_/B sky130_fd_sc_hd__or2_1
X_08905_ _08904_/X _08810_/B _08810_/Y VGND VGND VPWR VPWR _08905_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _10018_/A _10124_/A VGND VGND VPWR VPWR _08836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08767_ _09331_/B VGND VGND VPWR VPWR _10132_/A sky130_fd_sc_hd__clkbuf_2
X_08698_ _10008_/A VGND VGND VPWR VPWR _09478_/A sky130_fd_sc_hd__buf_1
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10660_ _11936_/A VGND VGND VPWR VPWR _13636_/A sky130_fd_sc_hd__buf_1
XFILLER_41_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09319_ _09531_/A _09737_/A VGND VGND VPWR VPWR _09353_/A sky130_fd_sc_hd__or2_1
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10591_ _09720_/A _09720_/B _09720_/Y VGND VGND VPWR VPWR _10592_/A sky130_fd_sc_hd__o21ai_1
X_12330_ _12240_/X _12329_/Y _12240_/X _12329_/Y VGND VGND VPWR VPWR _12590_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12261_ _12261_/A _12261_/B VGND VGND VPWR VPWR _12261_/X sky130_fd_sc_hd__and2_1
XFILLER_5_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11212_ _11087_/X _11211_/X _11087_/X _11211_/X VGND VGND VPWR VPWR _11213_/B sky130_fd_sc_hd__a2bb2o_1
X_14000_ _13994_/A _13994_/B _13994_/Y VGND VGND VPWR VPWR _14000_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12192_ _12256_/A _12256_/B VGND VGND VPWR VPWR _12192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11143_ _10082_/X _11142_/X _10082_/X _11142_/X VGND VGND VPWR VPWR _11144_/B sky130_fd_sc_hd__a2bb2o_1
X_15951_ _15942_/X _15949_/X _16020_/B VGND VGND VPWR VPWR _15951_/X sky130_fd_sc_hd__o21a_1
X_11074_ _14429_/A _11075_/B VGND VGND VPWR VPWR _11074_/X sky130_fd_sc_hd__or2_1
XFILLER_88_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15882_ _14231_/Y _15840_/A _14231_/Y _15840_/A VGND VGND VPWR VPWR _15886_/B sky130_fd_sc_hd__a2bb2o_1
X_14902_ _14815_/A _14815_/B _14815_/Y VGND VGND VPWR VPWR _14902_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10025_ _09492_/A _10128_/A _10050_/B _10024_/X VGND VGND VPWR VPWR _10025_/X sky130_fd_sc_hd__o22a_1
XFILLER_48_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14833_ _14833_/A _14833_/B VGND VGND VPWR VPWR _14833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14764_ _14833_/A _14833_/B VGND VGND VPWR VPWR _14764_/Y sky130_fd_sc_hd__nand2_1
X_11976_ _11976_/A _11976_/B VGND VGND VPWR VPWR _11976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14695_ _14736_/A _14736_/B VGND VGND VPWR VPWR _14784_/A sky130_fd_sc_hd__and2_1
X_13715_ _13715_/A _13778_/B VGND VGND VPWR VPWR _13715_/Y sky130_fd_sc_hd__nand2_1
X_10927_ _09436_/A _09436_/B _09436_/Y VGND VGND VPWR VPWR _10928_/A sky130_fd_sc_hd__o21ai_1
X_16434_ _16434_/A _16434_/B VGND VGND VPWR VPWR _16434_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13646_ _15044_/A _13506_/B _13506_/Y VGND VGND VPWR VPWR _13646_/Y sky130_fd_sc_hd__o21ai_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10858_ _09271_/A _10857_/A _09274_/A _10857_/Y _10929_/A VGND VGND VPWR VPWR _12061_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16365_ _16357_/X _16464_/Q _16358_/X _16407_/C _16361_/X VGND VGND VPWR VPWR _16464_/D
+ sky130_fd_sc_hd__o221a_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13577_ _12845_/A _13559_/B _13560_/Y _13576_/X VGND VGND VPWR VPWR _13577_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10789_ _09968_/Y _10788_/A _10079_/A _10788_/Y _10943_/A VGND VGND VPWR VPWR _12070_/A
+ sky130_fd_sc_hd__a221o_2
X_16296_ _16328_/A _16328_/B VGND VGND VPWR VPWR _16296_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12528_ _12527_/A _12527_/B _12527_/Y _12503_/X VGND VGND VPWR VPWR _12634_/B sky130_fd_sc_hd__o211a_1
X_15316_ _15275_/X _15315_/Y _15275_/X _15315_/Y VGND VGND VPWR VPWR _15337_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15247_ _15193_/A _15193_/B _15193_/Y VGND VGND VPWR VPWR _15247_/Y sky130_fd_sc_hd__o21ai_1
X_12459_ _15285_/A _12462_/B VGND VGND VPWR VPWR _12459_/X sky130_fd_sc_hd__and2_1
XFILLER_113_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15178_ _15178_/A _15178_/B VGND VGND VPWR VPWR _15178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14129_ _14060_/X _14128_/Y _14060_/X _14128_/Y VGND VGND VPWR VPWR _14132_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09670_ _09523_/X _09669_/X _09523_/X _09669_/X VGND VGND VPWR VPWR _10763_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_67_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08621_ _08717_/B VGND VGND VPWR VPWR _08623_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08552_ _09531_/A VGND VGND VPWR VPWR _09470_/B sky130_fd_sc_hd__inv_2
XFILLER_63_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08483_ _08276_/Y _08279_/B _08482_/X VGND VGND VPWR VPWR _08483_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09104_ _09407_/A _09104_/B VGND VGND VPWR VPWR _09104_/X sky130_fd_sc_hd__and2_1
XFILLER_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09035_ _09553_/B _09035_/B VGND VGND VPWR VPWR _09036_/B sky130_fd_sc_hd__or2_1
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09937_ _09937_/A _09937_/B VGND VGND VPWR VPWR _09937_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09868_ _09452_/Y _09867_/X _09470_/X VGND VGND VPWR VPWR _09868_/X sky130_fd_sc_hd__o21a_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09799_ _09799_/A _09799_/B VGND VGND VPWR VPWR _09834_/A sky130_fd_sc_hd__or2_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08819_ _08819_/A _10126_/A VGND VGND VPWR VPWR _08819_/Y sky130_fd_sc_hd__nor2_1
X_11830_ _13605_/A _11840_/B VGND VGND VPWR VPWR _11830_/Y sky130_fd_sc_hd__nor2_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11761_ _11760_/A _11760_/B _11760_/X _11753_/B VGND VGND VPWR VPWR _11806_/B sky130_fd_sc_hd__a22o_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10712_ _13068_/A VGND VGND VPWR VPWR _11976_/A sky130_fd_sc_hd__buf_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13500_ _13500_/A _13500_/B VGND VGND VPWR VPWR _13500_/Y sky130_fd_sc_hd__nand2_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14480_/A VGND VGND VPWR VPWR _15196_/A sky130_fd_sc_hd__buf_1
X_11692_ _11692_/A VGND VGND VPWR VPWR _11692_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13431_ _13427_/Y _13429_/Y _13430_/Y VGND VGND VPWR VPWR _13435_/B sky130_fd_sc_hd__o21ai_2
X_10643_ _10596_/Y _10641_/Y _10642_/Y VGND VGND VPWR VPWR _10644_/A sky130_fd_sc_hd__o21ai_2
X_16150_ _15718_/X _16150_/B VGND VGND VPWR VPWR _16150_/X sky130_fd_sc_hd__and2b_1
X_13362_ _13362_/A _13362_/B VGND VGND VPWR VPWR _13362_/X sky130_fd_sc_hd__or2_1
X_10574_ _10675_/A _11921_/A VGND VGND VPWR VPWR _10574_/Y sky130_fd_sc_hd__nor2_1
X_16081_ _16028_/X _16080_/X _16028_/X _16080_/X VGND VGND VPWR VPWR _16084_/B sky130_fd_sc_hd__a2bb2o_1
X_12313_ _12245_/X _12312_/Y _12245_/X _12312_/Y VGND VGND VPWR VPWR _12314_/B sky130_fd_sc_hd__a2bb2o_1
X_15101_ _12274_/X _15048_/X _12276_/B VGND VGND VPWR VPWR _15101_/X sky130_fd_sc_hd__o21a_1
Xrebuffer8 rebuffer9/X VGND VGND VPWR VPWR rebuffer8/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13293_ _13293_/A VGND VGND VPWR VPWR _13293_/Y sky130_fd_sc_hd__inv_2
X_15032_ _15032_/A _15032_/B VGND VGND VPWR VPWR _15032_/X sky130_fd_sc_hd__or2_1
X_12244_ _12220_/A _12220_/B _12220_/Y _12243_/X VGND VGND VPWR VPWR _12244_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12175_ _12174_/A _12174_/B _12174_/X _12089_/B VGND VGND VPWR VPWR _12268_/B sky130_fd_sc_hd__a22o_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11126_ _12944_/A VGND VGND VPWR VPWR _12189_/A sky130_fd_sc_hd__inv_2
XFILLER_122_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15934_ _15892_/A _15892_/B _15892_/Y VGND VGND VPWR VPWR _15934_/Y sky130_fd_sc_hd__o21ai_1
X_11057_ _13184_/A _10912_/B _10912_/Y VGND VGND VPWR VPWR _11057_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15865_ _15898_/A _15898_/B VGND VGND VPWR VPWR _15865_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10008_ _10008_/A _10008_/B VGND VGND VPWR VPWR _10008_/X sky130_fd_sc_hd__or2_1
X_14816_ _14815_/A _14815_/B _14046_/X _14815_/Y VGND VGND VPWR VPWR _14816_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15796_ _15792_/Y _16227_/A _15795_/Y VGND VGND VPWR VPWR _15800_/B sky130_fd_sc_hd__o21ai_1
XFILLER_64_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14747_ _15237_/A VGND VGND VPWR VPWR _14833_/A sky130_fd_sc_hd__buf_1
X_11959_ _11894_/X _11958_/Y _11894_/X _11958_/Y VGND VGND VPWR VPWR _11966_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14678_ _14669_/X _14677_/X _14669_/X _14677_/X VGND VGND VPWR VPWR _14680_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16417_ _16466_/Q VGND VGND VPWR VPWR _16437_/B sky130_fd_sc_hd__inv_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13629_ _15131_/A _13629_/B VGND VGND VPWR VPWR _13629_/Y sky130_fd_sc_hd__nand2_1
X_16348_ _16336_/A _16336_/B _16336_/Y VGND VGND VPWR VPWR _16348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16279_ _16273_/A _16338_/A _16273_/Y VGND VGND VPWR VPWR _16279_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09722_ _09723_/A _09723_/B VGND VGND VPWR VPWR _09722_/Y sky130_fd_sc_hd__nor2_1
X_09653_ _09615_/Y _09651_/X _09652_/Y VGND VGND VPWR VPWR _09653_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08604_ _09217_/B VGND VGND VPWR VPWR _08604_/Y sky130_fd_sc_hd__inv_2
X_09584_ _09557_/X _09583_/X _09557_/X _09583_/X VGND VGND VPWR VPWR _09662_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _08535_/A VGND VGND VPWR VPWR _08535_/Y sky130_fd_sc_hd__inv_2
X_08466_ _08465_/A _08239_/Y _08465_/Y _08239_/A _08441_/X VGND VGND VPWR VPWR _09146_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08397_ _08399_/B _08392_/A _08282_/A _08392_/Y _08663_/B VGND VGND VPWR VPWR _08398_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10290_ _13478_/A _10286_/B _10289_/X VGND VGND VPWR VPWR _10291_/B sky130_fd_sc_hd__o21ai_1
XFILLER_2_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09018_ _08778_/A _09014_/Y _09014_/Y _08558_/Y VGND VGND VPWR VPWR _09019_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13980_ _14836_/A _13980_/B VGND VGND VPWR VPWR _13980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12931_ _12904_/Y _12929_/X _12930_/Y VGND VGND VPWR VPWR _12931_/X sky130_fd_sc_hd__o21a_1
X_15650_ _15650_/A VGND VGND VPWR VPWR _15650_/Y sky130_fd_sc_hd__inv_2
X_12862_ _12793_/Y _12860_/X _12861_/Y VGND VGND VPWR VPWR _12862_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14601_ _14592_/X _14600_/X _14592_/X _14600_/X VGND VGND VPWR VPWR _14603_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11813_ _11813_/A _11813_/B VGND VGND VPWR VPWR _11814_/B sky130_fd_sc_hd__or2_1
X_15581_ _15700_/A _15581_/B VGND VGND VPWR VPWR _16051_/A sky130_fd_sc_hd__or2_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12793_ _13872_/A _12861_/B VGND VGND VPWR VPWR _12793_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14531_/A _14531_/B _14531_/Y VGND VGND VPWR VPWR _14532_/X sky130_fd_sc_hd__a21o_1
X_11744_ _11774_/A _11744_/B VGND VGND VPWR VPWR _11744_/X sky130_fd_sc_hd__or2_1
XFILLER_42_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11675_ _14143_/A _11567_/B _11567_/Y _11569_/A VGND VGND VPWR VPWR _12644_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14450_/Y _14461_/X _14462_/Y VGND VGND VPWR VPWR _14463_/X sky130_fd_sc_hd__o21a_1
XFILLER_41_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16202_ _16257_/A _16258_/B VGND VGND VPWR VPWR _16202_/Y sky130_fd_sc_hd__nor2_1
X_13414_ _13356_/X _13413_/X _13356_/X _13413_/X VGND VGND VPWR VPWR _13414_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10626_ _10626_/A _12920_/A VGND VGND VPWR VPWR _12043_/A sky130_fd_sc_hd__or2_1
XFILLER_127_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16133_ _16061_/X _16133_/B VGND VGND VPWR VPWR _16133_/X sky130_fd_sc_hd__and2b_1
X_14394_ _14311_/X _14392_/X _15590_/B VGND VGND VPWR VPWR _14394_/X sky130_fd_sc_hd__o21a_1
X_13345_ _13348_/A VGND VGND VPWR VPWR _15470_/A sky130_fd_sc_hd__buf_1
X_10557_ _10556_/Y _10453_/X _10464_/Y VGND VGND VPWR VPWR _10557_/X sky130_fd_sc_hd__o21a_1
X_16064_ _16121_/A _16121_/B VGND VGND VPWR VPWR _16138_/A sky130_fd_sc_hd__and2_1
X_13276_ _14724_/A _13276_/B VGND VGND VPWR VPWR _13276_/Y sky130_fd_sc_hd__nand2_1
X_10488_ _13624_/A _10531_/B VGND VGND VPWR VPWR _10488_/Y sky130_fd_sc_hd__nor2_1
X_12227_ _12227_/A _12141_/X VGND VGND VPWR VPWR _12227_/X sky130_fd_sc_hd__or2b_1
X_15015_ _11863_/Y _15002_/X _11863_/Y _15002_/X VGND VGND VPWR VPWR _15038_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12158_ _12157_/Y _12066_/X _12106_/Y VGND VGND VPWR VPWR _12158_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11109_ _12198_/A VGND VGND VPWR VPWR _11279_/A sky130_fd_sc_hd__inv_2
XFILLER_77_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12089_ _12089_/A _12089_/B VGND VGND VPWR VPWR _12089_/X sky130_fd_sc_hd__or2_1
X_15917_ _15907_/X _15916_/Y _15907_/X _15916_/Y VGND VGND VPWR VPWR _15970_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15848_ _14189_/A _15847_/X _12632_/X VGND VGND VPWR VPWR _15848_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15779_ _15777_/Y _15778_/Y _15777_/Y _15778_/Y VGND VGND VPWR VPWR _15785_/B sky130_fd_sc_hd__o2bb2a_1
X_08320_ _08318_/Y _08319_/A _08318_/A _08319_/Y _08304_/X VGND VGND VPWR VPWR _08543_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08251_ input3/X _08251_/B VGND VGND VPWR VPWR _08322_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09705_ _09705_/A VGND VGND VPWR VPWR _09720_/A sky130_fd_sc_hd__inv_2
XFILLER_114_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09636_ _09952_/A _09631_/B _09632_/Y _09635_/Y VGND VGND VPWR VPWR _09640_/B sky130_fd_sc_hd__o22a_1
XFILLER_82_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09567_ _09567_/A _09567_/B VGND VGND VPWR VPWR _09567_/X sky130_fd_sc_hd__or2_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08518_ _08701_/A _08518_/B VGND VGND VPWR VPWR _09525_/A sky130_fd_sc_hd__or2_2
X_09498_ _09498_/A _09498_/B VGND VGND VPWR VPWR _09498_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08449_ _08543_/A VGND VGND VPWR VPWR _10010_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11460_ _14131_/A _11365_/B _11365_/Y _12516_/A VGND VGND VPWR VPWR _12508_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10411_ _10411_/A VGND VGND VPWR VPWR _10411_/Y sky130_fd_sc_hd__inv_2
X_11391_ _08912_/X _11391_/B VGND VGND VPWR VPWR _11391_/X sky130_fd_sc_hd__and2b_1
XFILLER_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13130_ _13128_/Y _13129_/X _13128_/Y _13129_/X VGND VGND VPWR VPWR _13130_/X sky130_fd_sc_hd__o2bb2a_1
X_10342_ _13478_/A _10286_/B _10289_/A VGND VGND VPWR VPWR _10342_/X sky130_fd_sc_hd__o21ba_1
XFILLER_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13061_ _13026_/X _13060_/X _13026_/X _13060_/X VGND VGND VPWR VPWR _13117_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12012_ _12071_/A _12011_/Y _12071_/A _12011_/Y VGND VGND VPWR VPWR _12068_/B sky130_fd_sc_hd__a2bb2o_1
X_10273_ _10108_/Y _10272_/Y _10108_/A _10272_/A _10471_/A VGND VGND VPWR VPWR _11732_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15702_ _14403_/X _15701_/Y _14403_/X _15701_/Y VGND VGND VPWR VPWR _15825_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13963_ _13988_/A VGND VGND VPWR VPWR _14956_/A sky130_fd_sc_hd__buf_1
XFILLER_58_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13894_ _14663_/A _13857_/B _13857_/Y VGND VGND VPWR VPWR _13894_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12914_ _10425_/A _12834_/Y _10425_/A _12834_/Y VGND VGND VPWR VPWR _12915_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ _15633_/A VGND VGND VPWR VPWR _15633_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12845_ _12845_/A _12845_/B VGND VGND VPWR VPWR _12845_/Y sky130_fd_sc_hd__nand2_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15563_/Y _15486_/X _15433_/Y VGND VGND VPWR VPWR _15564_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12776_ _12776_/A _12776_/B VGND VGND VPWR VPWR _12776_/Y sky130_fd_sc_hd__nand2_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _15202_/A _14515_/B VGND VGND VPWR VPWR _14515_/X sky130_fd_sc_hd__or2_1
X_11727_ _11727_/A _11733_/A VGND VGND VPWR VPWR _11727_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15495_ _15443_/A _15443_/B _15443_/A _15443_/B VGND VGND VPWR VPWR _15495_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11658_ _11655_/X _11658_/B VGND VGND VPWR VPWR _11658_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_80_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14446_ _14433_/X _14445_/X _14433_/X _14445_/X VGND VGND VPWR VPWR _14464_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14377_ _14377_/A _14377_/B VGND VGND VPWR VPWR _14377_/Y sky130_fd_sc_hd__nand2_1
X_11589_ _09667_/Y _11588_/Y _09667_/Y _11588_/Y VGND VGND VPWR VPWR _11590_/B sky130_fd_sc_hd__o2bb2a_1
X_10609_ _09407_/A _09709_/B _09709_/Y VGND VGND VPWR VPWR _10610_/A sky130_fd_sc_hd__o21ai_1
XFILLER_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16116_ _16119_/A _16119_/B VGND VGND VPWR VPWR _16116_/Y sky130_fd_sc_hd__nor2_1
X_13328_ _13362_/A _13362_/B VGND VGND VPWR VPWR _13390_/A sky130_fd_sc_hd__and2_1
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16047_ _16001_/Y _16045_/X _16046_/Y VGND VGND VPWR VPWR _16051_/B sky130_fd_sc_hd__o21ai_2
X_13259_ _13187_/X _13258_/Y _13187_/X _13258_/Y VGND VGND VPWR VPWR _13279_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09421_ _09421_/A _09421_/B VGND VGND VPWR VPWR _09421_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09352_ _09352_/A VGND VGND VPWR VPWR _09352_/Y sky130_fd_sc_hd__inv_2
X_08303_ _08303_/A VGND VGND VPWR VPWR _08304_/A sky130_fd_sc_hd__clkbuf_2
X_09283_ _09462_/B _09801_/A _09227_/X VGND VGND VPWR VPWR _09283_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08234_ input23/X VGND VGND VPWR VPWR _08235_/B sky130_fd_sc_hd__inv_4
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08998_ _12606_/B VGND VGND VPWR VPWR _11411_/B sky130_fd_sc_hd__inv_2
XFILLER_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10960_ _10081_/A _10958_/Y _09967_/Y _10958_/A _10959_/X VGND VGND VPWR VPWR _12080_/A
+ sky130_fd_sc_hd__o221a_1
X_10891_ _12039_/A VGND VGND VPWR VPWR _13824_/A sky130_fd_sc_hd__buf_1
XFILLER_71_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09619_ _09500_/A _09500_/B _09500_/Y VGND VGND VPWR VPWR _09619_/X sky130_fd_sc_hd__a21o_1
X_12630_ _12630_/A _12630_/B VGND VGND VPWR VPWR _12630_/X sky130_fd_sc_hd__or2_1
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12561_ _12561_/A VGND VGND VPWR VPWR _12561_/Y sky130_fd_sc_hd__inv_2
X_14300_ _13443_/A _13443_/B _13443_/Y VGND VGND VPWR VPWR _14300_/X sky130_fd_sc_hd__o21a_1
X_12492_ _13132_/A _12488_/B _12488_/Y VGND VGND VPWR VPWR _12492_/Y sky130_fd_sc_hd__o21ai_1
X_15280_ _14587_/A _15246_/B _15246_/Y _15279_/X VGND VGND VPWR VPWR _15280_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11512_ _09964_/X _11512_/B VGND VGND VPWR VPWR _11513_/B sky130_fd_sc_hd__and2b_1
X_14231_ _14231_/A _12618_/X VGND VGND VPWR VPWR _14231_/Y sky130_fd_sc_hd__nor2b_1
X_11443_ _15529_/A _11443_/B VGND VGND VPWR VPWR _11443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14162_ _12650_/Y _14162_/B VGND VGND VPWR VPWR _14162_/X sky130_fd_sc_hd__and2b_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13113_ _15252_/A _13113_/B VGND VGND VPWR VPWR _13113_/Y sky130_fd_sc_hd__nand2_1
X_11374_ _08975_/X _11373_/X _08975_/X _11373_/X VGND VGND VPWR VPWR _11375_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14093_ _15464_/A _14035_/B _14035_/A _14035_/B VGND VGND VPWR VPWR _14093_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_98_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10325_ _10325_/A _10325_/B VGND VGND VPWR VPWR _10325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13044_ _13796_/A VGND VGND VPWR VPWR _15237_/A sky130_fd_sc_hd__buf_1
X_10256_ _09312_/A _10254_/B _10255_/Y _10468_/A VGND VGND VPWR VPWR _10571_/A sky130_fd_sc_hd__o22a_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10187_ _10243_/B _10159_/B _10159_/Y _10685_/A VGND VGND VPWR VPWR _10822_/A sky130_fd_sc_hd__o2bb2a_1
X_14995_ _15752_/A VGND VGND VPWR VPWR _15728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13946_ _13920_/Y _13944_/X _13945_/Y VGND VGND VPWR VPWR _13946_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15616_ _15616_/A VGND VGND VPWR VPWR _15616_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_62_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13877_ _13865_/X _13876_/Y _13865_/X _13876_/Y VGND VGND VPWR VPWR _13980_/B sky130_fd_sc_hd__a2bb2o_1
X_12828_ _12837_/A VGND VGND VPWR VPWR _15087_/A sky130_fd_sc_hd__clkbuf_2
X_15547_ _15500_/X _15545_/X _15586_/B VGND VGND VPWR VPWR _15547_/X sky130_fd_sc_hd__o21a_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12707_/A _12707_/B _12707_/Y VGND VGND VPWR VPWR _12759_/X sky130_fd_sc_hd__a21o_1
X_15478_ _14802_/A _15461_/B _15461_/Y _15477_/X VGND VGND VPWR VPWR _15478_/X sky130_fd_sc_hd__a2bb2o_1
X_14429_ _14429_/A _14429_/B VGND VGND VPWR VPWR _14429_/X sky130_fd_sc_hd__and2_1
XFILLER_128_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09970_ _09970_/A VGND VGND VPWR VPWR _09970_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08921_ _08930_/A _09101_/A VGND VGND VPWR VPWR _08922_/B sky130_fd_sc_hd__or2_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08852_ _08852_/A _08856_/B VGND VGND VPWR VPWR _08913_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08783_ _10130_/A VGND VGND VPWR VPWR _08786_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09404_ _09404_/A VGND VGND VPWR VPWR _09404_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09335_ _08778_/A _08776_/Y _10041_/A _09334_/X VGND VGND VPWR VPWR _09335_/X sky130_fd_sc_hd__o22a_1
X_09266_ _09258_/X _08899_/Y _09258_/X _08899_/Y VGND VGND VPWR VPWR _10243_/A sky130_fd_sc_hd__o2bb2a_1
X_09197_ _09146_/X _09150_/S _08505_/B VGND VGND VPWR VPWR _09199_/A sky130_fd_sc_hd__o21ba_2
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11090_ _13905_/A _11090_/B VGND VGND VPWR VPWR _11090_/X sky130_fd_sc_hd__or2_1
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10110_ _10110_/A _10110_/B VGND VGND VPWR VPWR _10111_/A sky130_fd_sc_hd__or2_1
XFILLER_96_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10041_ _10041_/A _10041_/B VGND VGND VPWR VPWR _10041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14780_ _14780_/A _14738_/X VGND VGND VPWR VPWR _14780_/X sky130_fd_sc_hd__or2b_1
X_13800_ _13722_/X _13800_/B VGND VGND VPWR VPWR _13800_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11992_ _11992_/A _11992_/B VGND VGND VPWR VPWR _11992_/X sky130_fd_sc_hd__or2_1
XFILLER_84_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13731_ _13768_/A _13768_/B VGND VGND VPWR VPWR _13809_/A sky130_fd_sc_hd__and2_1
XFILLER_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10943_ _10943_/A VGND VGND VPWR VPWR _11593_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16450_ _16445_/X _16448_/X _16474_/Q _16449_/X VGND VGND VPWR VPWR _16450_/X sky130_fd_sc_hd__o22a_1
X_10874_ _12057_/A VGND VGND VPWR VPWR _10878_/A sky130_fd_sc_hd__inv_2
X_13662_ _13631_/A _13661_/Y _13631_/A _13661_/Y VGND VGND VPWR VPWR _13696_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16381_ _16316_/A _16316_/B _16316_/Y VGND VGND VPWR VPWR _16381_/Y sky130_fd_sc_hd__o21ai_1
X_12613_ _15509_/A _12320_/B _12321_/A VGND VGND VPWR VPWR _12614_/A sky130_fd_sc_hd__o21ai_1
X_15401_ _15465_/A _15399_/X _15400_/X VGND VGND VPWR VPWR _15401_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13593_ _13555_/A _13555_/B _13556_/A VGND VGND VPWR VPWR _13593_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12544_ _12543_/A _12543_/B _12543_/Y _12503_/A VGND VGND VPWR VPWR _12630_/B sky130_fd_sc_hd__o211a_1
XFILLER_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15332_ _15326_/Y _15330_/X _15331_/Y VGND VGND VPWR VPWR _15332_/X sky130_fd_sc_hd__o21a_1
X_15263_ _15218_/X _15262_/Y _15218_/X _15262_/Y VGND VGND VPWR VPWR _15264_/B sky130_fd_sc_hd__a2bb2o_1
X_12475_ _12434_/X _12474_/X _12434_/X _12474_/X VGND VGND VPWR VPWR _12475_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_6 _16361_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14214_ _12623_/X _14213_/X _12623_/X _14213_/X VGND VGND VPWR VPWR _14259_/B sky130_fd_sc_hd__a2bb2o_1
X_11426_ _11253_/X _11425_/Y _11253_/X _11425_/Y VGND VGND VPWR VPWR _12595_/A sky130_fd_sc_hd__a2bb2o_1
X_15194_ _15128_/A _15128_/B _15128_/Y VGND VGND VPWR VPWR _15194_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14145_ _14139_/X _14142_/Y _14407_/A _14144_/Y VGND VGND VPWR VPWR _14145_/X sky130_fd_sc_hd__o22a_1
X_11357_ _11263_/X _11356_/Y _11263_/X _11356_/Y VGND VGND VPWR VPWR _11358_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14076_ _14076_/A _14055_/X VGND VGND VPWR VPWR _14076_/X sky130_fd_sc_hd__or2b_1
X_10308_ _11762_/A _10369_/B _10307_/Y VGND VGND VPWR VPWR _10310_/A sky130_fd_sc_hd__o21ai_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13027_ _14523_/A _13027_/B VGND VGND VPWR VPWR _13027_/X sky130_fd_sc_hd__or2_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _11590_/A _11288_/B VGND VGND VPWR VPWR _13043_/A sky130_fd_sc_hd__or2_2
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10239_ _10239_/A _10239_/B VGND VGND VPWR VPWR _10239_/X sky130_fd_sc_hd__or2_1
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer18 rebuffer19/X VGND VGND VPWR VPWR rebuffer18/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14978_ _14971_/A _14938_/B _14938_/Y _14940_/X VGND VGND VPWR VPWR _14978_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer29 _08662_/A VGND VGND VPWR VPWR _08507_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13929_ _14645_/A _13839_/B _13839_/Y VGND VGND VPWR VPWR _13929_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09120_ _09418_/A _09123_/B VGND VGND VPWR VPWR _09120_/Y sky130_fd_sc_hd__nor2_1
X_09051_ _08712_/Y _09050_/Y _08734_/X VGND VGND VPWR VPWR _09052_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09953_ _08928_/A _09707_/Y _09627_/A _09681_/A VGND VGND VPWR VPWR _09955_/B sky130_fd_sc_hd__o22a_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _09884_/A _09884_/B VGND VGND VPWR VPWR _09885_/B sky130_fd_sc_hd__or2_1
X_08904_ _10015_/A VGND VGND VPWR VPWR _08904_/X sky130_fd_sc_hd__buf_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _09252_/B VGND VGND VPWR VPWR _10124_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08766_ _08765_/A _08742_/A _08765_/Y _08742_/Y VGND VGND VPWR VPWR _09331_/B sky130_fd_sc_hd__o22a_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08697_ _08697_/A VGND VGND VPWR VPWR _10008_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09318_ _08572_/A _09858_/A _09317_/Y _09243_/X VGND VGND VPWR VPWR _09318_/X sky130_fd_sc_hd__o22a_1
X_10590_ _11907_/A _10645_/B VGND VGND VPWR VPWR _10590_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09249_ _09249_/A _10127_/A VGND VGND VPWR VPWR _10073_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12260_ _12259_/Y _12166_/X _12189_/Y VGND VGND VPWR VPWR _12260_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11211_ _11211_/A _11088_/X VGND VGND VPWR VPWR _11211_/X sky130_fd_sc_hd__or2b_1
X_12191_ _12166_/X _12190_/Y _12166_/X _12190_/Y VGND VGND VPWR VPWR _12256_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11142_ _10043_/X _11142_/B VGND VGND VPWR VPWR _11142_/X sky130_fd_sc_hd__and2b_1
XFILLER_134_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15950_ _15950_/A _15950_/B VGND VGND VPWR VPWR _16020_/B sky130_fd_sc_hd__or2_1
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11073_ _11067_/A _11072_/X _11067_/A _11072_/X VGND VGND VPWR VPWR _11075_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15881_ _15881_/A VGND VGND VPWR VPWR _15886_/A sky130_fd_sc_hd__clkinvlp_2
X_14901_ _14901_/A _14906_/B VGND VGND VPWR VPWR _14901_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10024_ _09249_/A _08810_/B _10073_/B _10023_/X VGND VGND VPWR VPWR _10024_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14832_ _14832_/A VGND VGND VPWR VPWR _15353_/A sky130_fd_sc_hd__buf_1
XFILLER_49_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11975_ _11948_/Y _11973_/X _11974_/Y VGND VGND VPWR VPWR _11975_/X sky130_fd_sc_hd__o21a_1
X_14763_ _14748_/X _14762_/X _14748_/X _14762_/X VGND VGND VPWR VPWR _14833_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10926_ _11013_/A _10923_/X _10925_/X VGND VGND VPWR VPWR _10926_/X sky130_fd_sc_hd__o21a_1
X_14694_ _14658_/X _14693_/Y _14658_/X _14693_/Y VGND VGND VPWR VPWR _14736_/B sky130_fd_sc_hd__a2bb2o_1
X_13714_ _13709_/X _13713_/Y _13709_/X _13713_/Y VGND VGND VPWR VPWR _13778_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16433_ _16429_/B _16426_/A _16420_/X VGND VGND VPWR VPWR _16434_/B sky130_fd_sc_hd__a21bo_1
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13645_ _12853_/A _13583_/B _13644_/Y _13580_/X VGND VGND VPWR VPWR _13645_/X sky130_fd_sc_hd__o22a_1
X_10857_ _10857_/A VGND VGND VPWR VPWR _10857_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16364_ _16327_/X _16363_/Y _16327_/X _16363_/Y VGND VGND VPWR VPWR _16407_/C sky130_fd_sc_hd__a2bb2o_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _12843_/A _13563_/B _13564_/Y _13575_/X VGND VGND VPWR VPWR _13576_/X sky130_fd_sc_hd__o22a_1
X_10788_ _10788_/A VGND VGND VPWR VPWR _10788_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16295_ _16261_/X _16294_/Y _16261_/X _16294_/Y VGND VGND VPWR VPWR _16328_/B sky130_fd_sc_hd__o2bb2a_1
X_12527_ _12527_/A _12527_/B VGND VGND VPWR VPWR _12527_/Y sky130_fd_sc_hd__nand2_1
X_15315_ _14579_/A _15258_/B _15258_/Y VGND VGND VPWR VPWR _15315_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15246_ _15246_/A _15246_/B VGND VGND VPWR VPWR _15246_/Y sky130_fd_sc_hd__nand2_1
X_12458_ _12455_/X _12482_/A _12455_/X _12482_/A VGND VGND VPWR VPWR _12462_/B sky130_fd_sc_hd__a2bb2o_1
X_11409_ _11409_/A VGND VGND VPWR VPWR _11409_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15177_ _15158_/X _15176_/Y _15158_/X _15176_/Y VGND VGND VPWR VPWR _15178_/B sky130_fd_sc_hd__a2bb2o_1
X_12389_ _12370_/X _12388_/X _12370_/X _12388_/X VGND VGND VPWR VPWR _12451_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14128_ _14011_/X _14128_/B VGND VGND VPWR VPWR _14128_/Y sky130_fd_sc_hd__nand2b_1
X_14059_ _14059_/A _14059_/B VGND VGND VPWR VPWR _14059_/X sky130_fd_sc_hd__or2_1
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08620_ _09457_/B VGND VGND VPWR VPWR _08717_/B sky130_fd_sc_hd__inv_2
XFILLER_82_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08551_ _08589_/A _08551_/B VGND VGND VPWR VPWR _09531_/A sky130_fd_sc_hd__or2_2
XFILLER_62_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08482_ _08276_/Y _08279_/B _08481_/Y VGND VGND VPWR VPWR _08482_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09103_ _09101_/A _08677_/B _08664_/X _09102_/Y VGND VGND VPWR VPWR _09104_/B sky130_fd_sc_hd__o22a_1
XFILLER_129_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09034_ _09551_/B _09034_/B VGND VGND VPWR VPWR _09035_/B sky130_fd_sc_hd__or2_1
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09936_ _08703_/A _09873_/A _08704_/B VGND VGND VPWR VPWR _09936_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09867_ _08893_/X _08572_/A _09453_/Y _09866_/X VGND VGND VPWR VPWR _09867_/X sky130_fd_sc_hd__o22a_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08818_ _09250_/B VGND VGND VPWR VPWR _10126_/A sky130_fd_sc_hd__clkbuf_2
X_09798_ _09700_/Y _09727_/A _09700_/A _09727_/Y _10943_/A VGND VGND VPWR VPWR _11910_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08749_ _08749_/A VGND VGND VPWR VPWR _08749_/Y sky130_fd_sc_hd__inv_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11760_ _11760_/A _11760_/B VGND VGND VPWR VPWR _11760_/X sky130_fd_sc_hd__or2_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10711_ _10933_/A _10711_/B VGND VGND VPWR VPWR _13068_/A sky130_fd_sc_hd__or2_2
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11685_/X _11690_/X _11685_/X _11690_/X VGND VGND VPWR VPWR _11691_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13430_ _14105_/A _13430_/B VGND VGND VPWR VPWR _13430_/Y sky130_fd_sc_hd__nand2_1
X_10642_ _11904_/A _10642_/B VGND VGND VPWR VPWR _10642_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13361_ _13331_/A _13331_/B _13331_/X _13360_/X VGND VGND VPWR VPWR _13361_/X sky130_fd_sc_hd__o22a_1
X_10573_ _11921_/A VGND VGND VPWR VPWR _12695_/A sky130_fd_sc_hd__buf_1
X_16080_ _16027_/A _16027_/B _16027_/Y VGND VGND VPWR VPWR _16080_/X sky130_fd_sc_hd__o21a_1
X_12312_ _14020_/A _12214_/B _12214_/Y VGND VGND VPWR VPWR _12312_/Y sky130_fd_sc_hd__o21ai_1
X_13292_ _13240_/Y _13290_/Y _13291_/Y VGND VGND VPWR VPWR _13293_/A sky130_fd_sc_hd__o21ai_2
X_15100_ _15047_/X _15050_/X _15052_/B VGND VGND VPWR VPWR _15100_/X sky130_fd_sc_hd__o21a_1
Xrebuffer9 rebuffer9/A VGND VGND VPWR VPWR rebuffer9/X sky130_fd_sc_hd__dlygate4sd1_1
X_12243_ _14028_/A _12223_/B _12223_/Y _12242_/X VGND VGND VPWR VPWR _12243_/X sky130_fd_sc_hd__a2bb2o_1
X_15031_ _15079_/A _15029_/X _15030_/X VGND VGND VPWR VPWR _15031_/X sky130_fd_sc_hd__o21a_1
X_12174_ _12174_/A _12174_/B VGND VGND VPWR VPWR _12174_/X sky130_fd_sc_hd__or2_1
XFILLER_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11125_ _09919_/Y _11124_/X _09918_/X _09921_/B _10794_/X VGND VGND VPWR VPWR _12944_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_1_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15933_ _15956_/A _15956_/B VGND VGND VPWR VPWR _15933_/X sky130_fd_sc_hd__and2_1
XFILLER_110_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11056_ _15084_/A VGND VGND VPWR VPWR _12139_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10007_ _08704_/B _09792_/A _09146_/X _09793_/B VGND VGND VPWR VPWR _10007_/X sky130_fd_sc_hd__a22o_1
X_15864_ _14195_/X _15846_/X _14195_/X _15846_/X VGND VGND VPWR VPWR _15898_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15795_ _16094_/A _15795_/B VGND VGND VPWR VPWR _15795_/Y sky130_fd_sc_hd__nand2_1
X_14815_ _14815_/A _14815_/B VGND VGND VPWR VPWR _14815_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14746_ _14665_/X _14745_/Y _14683_/Y VGND VGND VPWR VPWR _14746_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11958_ _11895_/A _11895_/B _11895_/Y VGND VGND VPWR VPWR _11958_/Y sky130_fd_sc_hd__o21ai_1
X_10909_ _10909_/A VGND VGND VPWR VPWR _11067_/A sky130_fd_sc_hd__inv_2
X_11889_ _11889_/A _12043_/A VGND VGND VPWR VPWR _11961_/A sky130_fd_sc_hd__or2_1
X_14677_ _14676_/A _14676_/B _14676_/Y VGND VGND VPWR VPWR _14677_/X sky130_fd_sc_hd__a21o_1
X_16416_ _16467_/Q VGND VGND VPWR VPWR _16416_/Y sky130_fd_sc_hd__inv_2
X_13628_ _13628_/A VGND VGND VPWR VPWR _15131_/A sky130_fd_sc_hd__buf_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16347_ _08230_/X _16469_/Q _08233_/X _16392_/B _16343_/X VGND VGND VPWR VPWR _16469_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_118_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13559_ _13559_/A _13559_/B VGND VGND VPWR VPWR _13560_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16278_ _16276_/X _16278_/B VGND VGND VPWR VPWR _16278_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_133_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15229_ _15178_/A _15178_/B _15178_/Y _15228_/X VGND VGND VPWR VPWR _15229_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_114_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09721_ _09971_/A _09719_/Y _09720_/Y VGND VGND VPWR VPWR _09723_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09652_ _09978_/A _09652_/B VGND VGND VPWR VPWR _09652_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08603_ _09217_/A VGND VGND VPWR VPWR _10015_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09583_ _08690_/A _09017_/A _09530_/A VGND VGND VPWR VPWR _09583_/X sky130_fd_sc_hd__o21a_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ _09743_/A _08567_/B VGND VGND VPWR VPWR _08535_/A sky130_fd_sc_hd__or2_1
XFILLER_82_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08465_ _08465_/A VGND VGND VPWR VPWR _08465_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08396_ _09232_/A VGND VGND VPWR VPWR _08852_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09017_ _09017_/A VGND VGND VPWR VPWR _09529_/B sky130_fd_sc_hd__inv_2
XFILLER_124_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09919_ _09740_/A _09914_/Y _09861_/B VGND VGND VPWR VPWR _09919_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12930_ _12930_/A _12930_/B VGND VGND VPWR VPWR _12930_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12861_ _13872_/A _12861_/B VGND VGND VPWR VPWR _12861_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14600_ _14599_/A _14599_/B _14599_/Y VGND VGND VPWR VPWR _14600_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11812_ _11813_/A _11813_/B VGND VGND VPWR VPWR _11812_/X sky130_fd_sc_hd__and2_1
XFILLER_37_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15580_ _15547_/X _15579_/X _15547_/X _15579_/X VGND VGND VPWR VPWR _15581_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12785_/X _12791_/Y _12785_/X _12791_/Y VGND VGND VPWR VPWR _12861_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14531_/A _14531_/B VGND VGND VPWR VPWR _14531_/Y sky130_fd_sc_hd__nor2_1
X_11743_ _11779_/A _11731_/B _11731_/X _11742_/Y VGND VGND VPWR VPWR _11744_/B sky130_fd_sc_hd__a22o_1
XFILLER_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11674_ _15554_/A _11676_/B VGND VGND VPWR VPWR _11674_/X sky130_fd_sc_hd__and2_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14462_/A _14462_/B VGND VGND VPWR VPWR _14462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16201_ _16205_/A _16201_/B VGND VGND VPWR VPWR _16258_/B sky130_fd_sc_hd__or2_1
X_13413_ _15467_/A _13344_/B _13344_/Y VGND VGND VPWR VPWR _13413_/X sky130_fd_sc_hd__a21o_1
X_10625_ _10625_/A _12917_/A _10625_/C VGND VGND VPWR VPWR _12920_/A sky130_fd_sc_hd__and3_1
XFILLER_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16132_ _16189_/A VGND VGND VPWR VPWR _16388_/A sky130_fd_sc_hd__buf_1
X_14393_ _15964_/A _14393_/B VGND VGND VPWR VPWR _15590_/B sky130_fd_sc_hd__or2_1
XFILLER_127_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13344_ _13344_/A _13344_/B VGND VGND VPWR VPWR _13344_/Y sky130_fd_sc_hd__nor2_1
X_10556_ _11857_/A _10556_/B VGND VGND VPWR VPWR _10556_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16063_ _16052_/Y _16062_/Y _16052_/Y _16062_/Y VGND VGND VPWR VPWR _16121_/B sky130_fd_sc_hd__o2bb2a_1
X_13275_ _13268_/Y _13273_/X _13274_/Y VGND VGND VPWR VPWR _13275_/X sky130_fd_sc_hd__o21a_1
X_10487_ _10434_/X _10486_/X _10434_/X _10486_/X VGND VGND VPWR VPWR _10531_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12226_ _14032_/A _12226_/B VGND VGND VPWR VPWR _12226_/Y sky130_fd_sc_hd__nand2_1
X_15014_ _15040_/A _15040_/B VGND VGND VPWR VPWR _15064_/A sky130_fd_sc_hd__and2_1
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12157_ _13200_/A _12157_/B VGND VGND VPWR VPWR _12157_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11108_ _11107_/A _11106_/Y _11107_/Y _11106_/A _11586_/A VGND VGND VPWR VPWR _12198_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12088_ _12089_/A _12089_/B VGND VGND VPWR VPWR _12090_/A sky130_fd_sc_hd__and2_1
X_15916_ _15908_/A _15908_/B _15908_/Y VGND VGND VPWR VPWR _15916_/Y sky130_fd_sc_hd__o21ai_1
X_11039_ _10878_/A _10878_/B _10878_/A _10878_/B VGND VGND VPWR VPWR _11039_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15847_ _14195_/A _15846_/X _12630_/X VGND VGND VPWR VPWR _15847_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15778_ _15778_/A _15664_/X VGND VGND VPWR VPWR _15778_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_52_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14729_ _14800_/A _14727_/X _14728_/X VGND VGND VPWR VPWR _14729_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08250_ input19/X VGND VGND VPWR VPWR _08251_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_33_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09704_ _09692_/A _09692_/B _09695_/A VGND VGND VPWR VPWR _09971_/A sky130_fd_sc_hd__a21bo_1
XFILLER_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09635_ _09635_/A VGND VGND VPWR VPWR _09635_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09566_ _09999_/A VGND VGND VPWR VPWR _09569_/A sky130_fd_sc_hd__buf_1
X_08517_ _08516_/A _08313_/Y _08516_/Y _08313_/A VGND VGND VPWR VPWR _08518_/B sky130_fd_sc_hd__o22a_1
X_09497_ _08823_/X _09464_/X _08823_/X _09464_/X VGND VGND VPWR VPWR _09498_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08448_ _08447_/A _08318_/Y _08447_/Y _08318_/A _08441_/X VGND VGND VPWR VPWR _08543_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10410_ _09297_/A _09297_/B _09298_/A VGND VGND VPWR VPWR _10411_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08379_ _08298_/X _08378_/X _08298_/A _08378_/X VGND VGND VPWR VPWR _08662_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11390_ _14107_/A VGND VGND VPWR VPWR _12351_/A sky130_fd_sc_hd__inv_2
X_10341_ _11718_/A VGND VGND VPWR VPWR _12832_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13060_ _13060_/A _13027_/X VGND VGND VPWR VPWR _13060_/X sky130_fd_sc_hd__or2b_1
X_10272_ _10272_/A VGND VGND VPWR VPWR _10272_/Y sky130_fd_sc_hd__inv_2
X_12011_ _13700_/A _12070_/B _12010_/Y VGND VGND VPWR VPWR _12011_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13962_ _13888_/Y _13960_/X _13961_/Y VGND VGND VPWR VPWR _13962_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15701_ _15982_/A _14404_/B _14404_/Y VGND VGND VPWR VPWR _15701_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12913_ _13609_/A VGND VGND VPWR VPWR _13005_/A sky130_fd_sc_hd__buf_1
X_13893_ _13893_/A VGND VGND VPWR VPWR _15416_/A sky130_fd_sc_hd__buf_1
XFILLER_74_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ _15632_/A VGND VGND VPWR VPWR _15632_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12844_ _12820_/Y _12842_/X _12843_/Y VGND VGND VPWR VPWR _12844_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15563_/A _15563_/B VGND VGND VPWR VPWR _15563_/Y sky130_fd_sc_hd__nor2_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12775_ _12745_/Y _12773_/X _12774_/Y VGND VGND VPWR VPWR _12775_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14556_/A _14512_/X _14513_/X VGND VGND VPWR VPWR _14514_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11726_ _12705_/A _11736_/B _12705_/A _11736_/B VGND VGND VPWR VPWR _11733_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15494_ _15550_/A _15550_/B VGND VGND VPWR VPWR _15494_/X sky130_fd_sc_hd__and2_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11657_ _13988_/A _11657_/B VGND VGND VPWR VPWR _11658_/B sky130_fd_sc_hd__or2_1
X_14445_ _14422_/A _14422_/B _14422_/Y VGND VGND VPWR VPWR _14445_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14376_ _15662_/B _14374_/Y _15661_/A VGND VGND VPWR VPWR _14376_/X sky130_fd_sc_hd__o21a_1
X_10608_ _11885_/A _10635_/B VGND VGND VPWR VPWR _10608_/Y sky130_fd_sc_hd__nor2_1
X_11588_ _09569_/A _09569_/B _09569_/Y VGND VGND VPWR VPWR _11588_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_128_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16115_ _16067_/X _16113_/X _16155_/B VGND VGND VPWR VPWR _16119_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13327_ _13290_/A _13326_/Y _13290_/A _13326_/Y VGND VGND VPWR VPWR _13362_/B sky130_fd_sc_hd__a2bb2o_1
X_10539_ _11848_/A VGND VGND VPWR VPWR _13555_/A sky130_fd_sc_hd__buf_1
XFILLER_6_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16046_ _16046_/A _16046_/B VGND VGND VPWR VPWR _16046_/Y sky130_fd_sc_hd__nand2_1
X_13258_ _13188_/A _13188_/B _13188_/Y VGND VGND VPWR VPWR _13258_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12209_ _12209_/A _12153_/X VGND VGND VPWR VPWR _12209_/X sky130_fd_sc_hd__or2b_1
X_13189_ _13171_/Y _13187_/X _13188_/Y VGND VGND VPWR VPWR _13189_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09420_ _09421_/A _09421_/B VGND VGND VPWR VPWR _09420_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09351_ _09529_/A _09740_/A VGND VGND VPWR VPWR _09352_/A sky130_fd_sc_hd__or2_1
X_09282_ _10250_/A VGND VGND VPWR VPWR _10252_/A sky130_fd_sc_hd__buf_1
X_08302_ _08663_/B VGND VGND VPWR VPWR _08303_/A sky130_fd_sc_hd__clkbuf_2
X_08233_ _08233_/A VGND VGND VPWR VPWR _08233_/X sky130_fd_sc_hd__buf_1
XFILLER_100_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08997_ _08997_/A VGND VGND VPWR VPWR _12606_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10890_ _12053_/A VGND VGND VPWR VPWR _12039_/A sky130_fd_sc_hd__buf_1
XFILLER_83_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09618_ _09974_/A VGND VGND VPWR VPWR _09975_/A sky130_fd_sc_hd__buf_1
XFILLER_71_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09549_ _09549_/A _09549_/B VGND VGND VPWR VPWR _09613_/B sky130_fd_sc_hd__and2_1
XFILLER_71_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12560_ _12556_/Y _12559_/Y _12556_/A _12559_/A _11710_/A VGND VGND VPWR VPWR _12626_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12491_ _12481_/Y _12490_/X _12481_/Y _12490_/X VGND VGND VPWR VPWR _12491_/X sky130_fd_sc_hd__a2bb2o_1
X_11511_ _13500_/A _11510_/B _11510_/X _11307_/X VGND VGND VPWR VPWR _11511_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14230_ _14230_/A _14230_/B VGND VGND VPWR VPWR _15881_/A sky130_fd_sc_hd__or2_1
X_11442_ _13395_/A VGND VGND VPWR VPWR _15529_/A sky130_fd_sc_hd__buf_1
X_14161_ _14281_/A _14161_/B VGND VGND VPWR VPWR _15974_/A sky130_fd_sc_hd__or2_1
XFILLER_109_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11373_ _08896_/X _11373_/B VGND VGND VPWR VPWR _11373_/X sky130_fd_sc_hd__and2b_1
XFILLER_125_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13112_ _13077_/Y _13110_/X _13111_/Y VGND VGND VPWR VPWR _13112_/X sky130_fd_sc_hd__o21a_1
X_10324_ _10324_/A VGND VGND VPWR VPWR _13527_/A sky130_fd_sc_hd__buf_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14092_ _14092_/A _14095_/B VGND VGND VPWR VPWR _14092_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13043_ _13043_/A VGND VGND VPWR VPWR _13796_/A sky130_fd_sc_hd__inv_2
X_10255_ _10255_/A VGND VGND VPWR VPWR _10255_/Y sky130_fd_sc_hd__inv_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10186_ _10244_/B _10163_/B _10163_/Y _10564_/A VGND VGND VPWR VPWR _10685_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_94_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14994_ _15766_/A VGND VGND VPWR VPWR _15752_/A sky130_fd_sc_hd__buf_6
X_13945_ _15404_/A _13945_/B VGND VGND VPWR VPWR _13945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13876_ _15110_/A _13974_/B _13875_/Y VGND VGND VPWR VPWR _13876_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15615_ _14914_/A _15534_/B _15534_/Y VGND VGND VPWR VPWR _15617_/A sky130_fd_sc_hd__o21ai_1
X_12827_ _12827_/A VGND VGND VPWR VPWR _12837_/A sky130_fd_sc_hd__inv_2
XFILLER_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15546_ _15546_/A _15546_/B VGND VGND VPWR VPWR _15586_/B sky130_fd_sc_hd__or2_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _15028_/A VGND VGND VPWR VPWR _12764_/A sky130_fd_sc_hd__inv_2
XFILLER_42_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11709_ _11709_/A VGND VGND VPWR VPWR _11710_/A sky130_fd_sc_hd__clkbuf_2
X_15477_ _14806_/A _15464_/B _15464_/Y _15476_/X VGND VGND VPWR VPWR _15477_/X sky130_fd_sc_hd__a2bb2o_1
X_12689_ _12689_/A _12689_/B VGND VGND VPWR VPWR _12689_/Y sky130_fd_sc_hd__nor2_1
X_14428_ _14428_/A _14428_/B VGND VGND VPWR VPWR _14428_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14359_ _15948_/A VGND VGND VPWR VPWR _14377_/B sky130_fd_sc_hd__inv_2
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16029_ _16027_/A _16027_/B _16027_/Y _16028_/X VGND VGND VPWR VPWR _16029_/X sky130_fd_sc_hd__a2bb2o_1
X_08920_ _09541_/A _09066_/A _09234_/A _09817_/B VGND VGND VPWR VPWR _09101_/A sky130_fd_sc_hd__o22a_2
X_08851_ _09677_/A VGND VGND VPWR VPWR _08916_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08782_ _08781_/A _08736_/A _08781_/Y _08736_/Y VGND VGND VPWR VPWR _10130_/A sky130_fd_sc_hd__o22a_1
XFILLER_84_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09403_ _09404_/A VGND VGND VPWR VPWR _09403_/X sky130_fd_sc_hd__clkbuf_2
X_09334_ _09470_/A _08784_/Y _10044_/A _09324_/X VGND VGND VPWR VPWR _09334_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09265_ _09265_/A VGND VGND VPWR VPWR _09268_/A sky130_fd_sc_hd__inv_2
XFILLER_21_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09196_ _09198_/A VGND VGND VPWR VPWR _09196_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10040_ _10085_/A _10085_/B VGND VGND VPWR VPWR _10040_/X sky130_fd_sc_hd__and2_1
XFILLER_102_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11991_ _12077_/A VGND VGND VPWR VPWR _12778_/A sky130_fd_sc_hd__buf_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13730_ _13697_/X _13729_/X _13697_/X _13729_/X VGND VGND VPWR VPWR _13768_/B sky130_fd_sc_hd__a2bb2o_1
X_10942_ _10942_/A VGND VGND VPWR VPWR _10942_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15400_ _15400_/A _15400_/B VGND VGND VPWR VPWR _15400_/X sky130_fd_sc_hd__or2_1
XFILLER_71_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13661_ _15128_/A _13633_/B _13633_/Y VGND VGND VPWR VPWR _13661_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10873_ _09946_/A _10872_/A _09946_/Y _10872_/Y _09445_/A VGND VGND VPWR VPWR _12057_/A
+ sky130_fd_sc_hd__a221o_2
X_16380_ _08230_/A _16459_/Q _08233_/A _16396_/A _16343_/A VGND VGND VPWR VPWR _16459_/D
+ sky130_fd_sc_hd__o221a_2
X_12612_ _14081_/A VGND VGND VPWR VPWR _15509_/A sky130_fd_sc_hd__buf_1
X_13592_ _13632_/A _13633_/B VGND VGND VPWR VPWR _13592_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12543_ _12543_/A _12543_/B VGND VGND VPWR VPWR _12543_/Y sky130_fd_sc_hd__nand2_1
X_15331_ _15331_/A _15331_/B VGND VGND VPWR VPWR _15331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15262_ _15208_/A _15208_/B _15208_/Y VGND VGND VPWR VPWR _15262_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14213_ _14213_/A _12624_/X VGND VGND VPWR VPWR _14213_/X sky130_fd_sc_hd__or2b_1
X_12474_ _12444_/Y _12473_/X _12444_/Y _12473_/X VGND VGND VPWR VPWR _12474_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 _16361_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11425_ _13348_/A _11244_/B _11244_/Y VGND VGND VPWR VPWR _11425_/Y sky130_fd_sc_hd__o21ai_1
X_15193_ _15193_/A _15193_/B VGND VGND VPWR VPWR _15193_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14144_ _14144_/A VGND VGND VPWR VPWR _14144_/Y sky130_fd_sc_hd__inv_2
X_11356_ _14063_/A _11355_/B _11355_/Y VGND VGND VPWR VPWR _11356_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14075_ _13977_/X _13981_/X _13979_/B VGND VGND VPWR VPWR _14075_/Y sky130_fd_sc_hd__o21ai_1
X_10307_ _11762_/A _10369_/B VGND VGND VPWR VPWR _10307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13026_ _13065_/A _13024_/X _13025_/X VGND VGND VPWR VPWR _13026_/X sky130_fd_sc_hd__o21a_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _09663_/X _11286_/X _09663_/X _11286_/X VGND VGND VPWR VPWR _11288_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10238_ _10238_/A _10238_/B VGND VGND VPWR VPWR _10238_/X sky130_fd_sc_hd__or2_1
XFILLER_67_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10169_ _10125_/A _10125_/B _10126_/B VGND VGND VPWR VPWR _10170_/B sky130_fd_sc_hd__a21bo_1
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14977_ _14976_/Y _14954_/X _14951_/Y VGND VGND VPWR VPWR _14977_/Y sky130_fd_sc_hd__o21ai_1
X_13928_ _15400_/A _13941_/B VGND VGND VPWR VPWR _13928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer19 rebuffer20/X VGND VGND VPWR VPWR rebuffer19/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_74_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13859_ _14744_/A _13859_/B VGND VGND VPWR VPWR _13859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15529_ _15529_/A _15529_/B VGND VGND VPWR VPWR _15529_/Y sky130_fd_sc_hd__nand2_1
X_09050_ _09050_/A VGND VGND VPWR VPWR _09050_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09952_ _09952_/A VGND VGND VPWR VPWR _09955_/A sky130_fd_sc_hd__inv_2
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08903_ _08684_/X _08902_/X _08684_/X _08902_/X VGND VGND VPWR VPWR _08972_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09883_/A _09883_/B VGND VGND VPWR VPWR _09884_/B sky130_fd_sc_hd__or2_1
XFILLER_111_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08834_/A VGND VGND VPWR VPWR _09252_/B sky130_fd_sc_hd__inv_2
XFILLER_85_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08765_ _08765_/A VGND VGND VPWR VPWR _08765_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08696_ _08515_/X _08695_/Y _08515_/X _08695_/Y VGND VGND VPWR VPWR _08986_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09317_ _09317_/A VGND VGND VPWR VPWR _09317_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09248_ _09492_/A _09248_/B VGND VGND VPWR VPWR _10050_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09179_ _09179_/A VGND VGND VPWR VPWR _09179_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11210_ _14023_/A VGND VGND VPWR VPWR _14108_/A sky130_fd_sc_hd__buf_1
X_12190_ _13715_/A _12259_/B _12189_/Y VGND VGND VPWR VPWR _12190_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11141_ _11140_/Y _10967_/X _10978_/Y VGND VGND VPWR VPWR _11141_/X sky130_fd_sc_hd__o21a_1
XFILLER_134_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11072_ _12049_/A _10910_/B _10910_/Y VGND VGND VPWR VPWR _11072_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15880_ _15888_/A _15888_/B VGND VGND VPWR VPWR _15880_/Y sky130_fd_sc_hd__nor2_1
X_14900_ _14816_/X _14899_/X _14816_/X _14899_/X VGND VGND VPWR VPWR _14906_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10023_ _09456_/A _10126_/A _10069_/B _10022_/X VGND VGND VPWR VPWR _10023_/X sky130_fd_sc_hd__o22a_1
X_14831_ _14743_/X _14830_/Y _14767_/Y VGND VGND VPWR VPWR _14831_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11974_ _11974_/A _11974_/B VGND VGND VPWR VPWR _11974_/Y sky130_fd_sc_hd__nand2_1
X_14762_ _14762_/A _14761_/X VGND VGND VPWR VPWR _14762_/X sky130_fd_sc_hd__or2b_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14693_ _15345_/A _14659_/B _14659_/Y VGND VGND VPWR VPWR _14693_/Y sky130_fd_sc_hd__o21ai_1
X_10925_ _14610_/A _10925_/B VGND VGND VPWR VPWR _10925_/X sky130_fd_sc_hd__or2_1
XFILLER_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13713_ _13712_/A _13712_/B _13781_/A VGND VGND VPWR VPWR _13713_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16432_ _16445_/A _16431_/Y _16445_/A _16431_/Y VGND VGND VPWR VPWR _16432_/X sky130_fd_sc_hd__a2bb2o_1
X_13644_ _13644_/A VGND VGND VPWR VPWR _13644_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10856_ _09421_/A _09421_/B _09421_/Y VGND VGND VPWR VPWR _10857_/A sky130_fd_sc_hd__o21ai_1
X_16363_ _16328_/A _16328_/B _16328_/Y VGND VGND VPWR VPWR _16363_/Y sky130_fd_sc_hd__o21ai_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ _15339_/A _15339_/B VGND VGND VPWR VPWR _15378_/A sky130_fd_sc_hd__and2_1
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _12841_/A _13567_/B _13568_/Y _13574_/Y VGND VGND VPWR VPWR _13575_/X sky130_fd_sc_hd__o22a_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10787_ _09776_/A _09776_/B _09776_/Y VGND VGND VPWR VPWR _10788_/A sky130_fd_sc_hd__o21ai_1
X_16294_ _16262_/A _16328_/A _16262_/Y VGND VGND VPWR VPWR _16294_/Y sky130_fd_sc_hd__o21ai_1
X_12526_ _13441_/A _12308_/B _12308_/Y VGND VGND VPWR VPWR _12527_/B sky130_fd_sc_hd__o21a_1
X_15245_ _15224_/X _15244_/Y _15224_/X _15244_/Y VGND VGND VPWR VPWR _15246_/B sky130_fd_sc_hd__a2bb2o_1
X_12457_ _12456_/Y _12366_/X _12393_/Y VGND VGND VPWR VPWR _12482_/A sky130_fd_sc_hd__o21ai_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15176_ _15110_/A _15110_/B _15110_/Y VGND VGND VPWR VPWR _15176_/Y sky130_fd_sc_hd__o21ai_1
X_11408_ _08942_/A _08942_/B _08942_/Y VGND VGND VPWR VPWR _11409_/A sky130_fd_sc_hd__o21ai_1
XFILLER_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14127_ _14121_/X _14124_/Y _14872_/A _14126_/Y VGND VGND VPWR VPWR _14127_/X sky130_fd_sc_hd__o22a_1
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12388_ _13871_/A _12442_/B _13871_/A _12442_/B VGND VGND VPWR VPWR _12388_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11339_ _11305_/X _11338_/X _11305_/X _11338_/X VGND VGND VPWR VPWR _11500_/B sky130_fd_sc_hd__a2bb2o_1
X_14058_ _14116_/A _14056_/X _14057_/X VGND VGND VPWR VPWR _14058_/X sky130_fd_sc_hd__o21a_1
X_13009_ _13009_/A VGND VGND VPWR VPWR _13009_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08550_ _08549_/A _08328_/Y _08549_/Y _08328_/A VGND VGND VPWR VPWR _08551_/B sky130_fd_sc_hd__o22a_1
XFILLER_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08481_ input2/X input18/X VGND VGND VPWR VPWR _08481_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09102_ _10102_/B _10098_/B VGND VGND VPWR VPWR _09102_/Y sky130_fd_sc_hd__nor2_1
X_09033_ _09549_/B _09033_/B VGND VGND VPWR VPWR _09034_/B sky130_fd_sc_hd__or2_1
XFILLER_116_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09935_ _09864_/X _09933_/X _09934_/X VGND VGND VPWR VPWR _09935_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_131_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09866_ _09454_/Y _09865_/X _09467_/X VGND VGND VPWR VPWR _09866_/X sky130_fd_sc_hd__o21a_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08817_ _08817_/A VGND VGND VPWR VPWR _09250_/B sky130_fd_sc_hd__inv_2
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09797_ _09797_/A VGND VGND VPWR VPWR _10943_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08748_ _09340_/B VGND VGND VPWR VPWR _08748_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08679_ _08679_/A _08679_/B VGND VGND VPWR VPWR _08679_/X sky130_fd_sc_hd__and2_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10710_ _09653_/X _10709_/X _09653_/X _10709_/X VGND VGND VPWR VPWR _10711_/B sky130_fd_sc_hd__a2bb2oi_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11687_/X _11689_/X _11687_/X _11689_/X VGND VGND VPWR VPWR _11690_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10641_ _10641_/A VGND VGND VPWR VPWR _10641_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13360_ _13334_/A _13334_/B _13334_/X _13359_/X VGND VGND VPWR VPWR _13360_/X sky130_fd_sc_hd__o22a_1
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10572_ _10571_/A _10571_/B _10571_/Y _10984_/A VGND VGND VPWR VPWR _11921_/A sky130_fd_sc_hd__o211a_1
XFILLER_22_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12311_ _12311_/A _12311_/B VGND VGND VPWR VPWR _12311_/Y sky130_fd_sc_hd__nand2_1
X_13291_ _14734_/A _13291_/B VGND VGND VPWR VPWR _13291_/Y sky130_fd_sc_hd__nand2_1
X_12242_ _14032_/A _12226_/B _12226_/Y _12241_/X VGND VGND VPWR VPWR _12242_/X sky130_fd_sc_hd__a2bb2o_1
X_15030_ _15030_/A _15030_/B VGND VGND VPWR VPWR _15030_/X sky130_fd_sc_hd__or2_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12173_ _12263_/A VGND VGND VPWR VPWR _12782_/A sky130_fd_sc_hd__buf_1
XFILLER_122_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11124_ _09918_/A _09918_/B _09918_/X VGND VGND VPWR VPWR _11124_/X sky130_fd_sc_hd__o21ba_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15932_ _15893_/X _15931_/Y _15893_/X _15931_/Y VGND VGND VPWR VPWR _15956_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11055_ _12826_/A VGND VGND VPWR VPWR _15084_/A sky130_fd_sc_hd__buf_1
XFILLER_1_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10006_ _11713_/A VGND VGND VPWR VPWR _13524_/A sky130_fd_sc_hd__buf_1
XFILLER_49_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15863_ _15863_/A VGND VGND VPWR VPWR _15898_/A sky130_fd_sc_hd__inv_2
XFILLER_67_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15794_ _15668_/Y _15793_/Y _15668_/Y _15793_/Y VGND VGND VPWR VPWR _16227_/A sky130_fd_sc_hd__a2bb2o_1
X_14814_ _13936_/X _14813_/Y _13936_/X _14813_/Y VGND VGND VPWR VPWR _14815_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14745_ _14745_/A _14745_/B VGND VGND VPWR VPWR _14745_/Y sky130_fd_sc_hd__nor2_1
X_11957_ _13088_/A _11968_/B VGND VGND VPWR VPWR _11957_/Y sky130_fd_sc_hd__nor2_1
X_10908_ _15212_/B _12043_/B VGND VGND VPWR VPWR _10909_/A sky130_fd_sc_hd__or2_1
X_16415_ _16415_/A VGND VGND VPWR VPWR _16415_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11888_ _11888_/A _11895_/B VGND VGND VPWR VPWR _11888_/Y sky130_fd_sc_hd__nor2_1
X_14676_ _14676_/A _14676_/B VGND VGND VPWR VPWR _14676_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13627_ _13627_/A VGND VGND VPWR VPWR _13627_/Y sky130_fd_sc_hd__inv_2
X_10839_ _12007_/A _10946_/B VGND VGND VPWR VPWR _10839_/Y sky130_fd_sc_hd__nand2_1
X_16346_ _16337_/X _16345_/Y _16337_/X _16345_/Y VGND VGND VPWR VPWR _16392_/B sky130_fd_sc_hd__a2bb2o_1
X_13558_ _13533_/X _13557_/Y _13533_/X _13557_/Y VGND VGND VPWR VPWR _13559_/B sky130_fd_sc_hd__a2bb2o_1
X_16277_ _16277_/A _16277_/B VGND VGND VPWR VPWR _16278_/B sky130_fd_sc_hd__or2_1
X_12509_ _12508_/A _12508_/B _12508_/Y _11710_/X VGND VGND VPWR VPWR _12638_/A sky130_fd_sc_hd__o211a_1
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15228_ _15181_/A _15181_/B _15181_/Y _15227_/X VGND VGND VPWR VPWR _15228_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13489_ _11136_/Y _12089_/A _10987_/Y _13488_/X VGND VGND VPWR VPWR _13489_/X sky130_fd_sc_hd__o22a_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15159_ _15110_/A _15110_/B _15110_/Y _15158_/X VGND VGND VPWR VPWR _15159_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09720_ _09720_/A _09720_/B VGND VGND VPWR VPWR _09720_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09651_ _09647_/Y _10726_/A _09650_/Y VGND VGND VPWR VPWR _09651_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08602_ _09456_/B VGND VGND VPWR VPWR _09549_/A sky130_fd_sc_hd__buf_1
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09582_ _09992_/A VGND VGND VPWR VPWR _09993_/A sky130_fd_sc_hd__buf_1
XFILLER_36_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08533_ _09861_/A VGND VGND VPWR VPWR _09743_/A sky130_fd_sc_hd__inv_2
XFILLER_63_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08464_ _08464_/A VGND VGND VPWR VPWR _08464_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08395_ _08395_/A VGND VGND VPWR VPWR _09232_/A sky130_fd_sc_hd__inv_2
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09016_ _08770_/A _09015_/X _09015_/X _08546_/Y VGND VGND VPWR VPWR _09017_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09918_ _09918_/A _09918_/B VGND VGND VPWR VPWR _09918_/X sky130_fd_sc_hd__and2_1
XFILLER_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09849_ _09693_/A _09844_/Y _09803_/B VGND VGND VPWR VPWR _09849_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12860_ _12796_/Y _12858_/X _12859_/Y VGND VGND VPWR VPWR _12860_/X sky130_fd_sc_hd__o21a_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11811_ _10466_/A _11810_/A _10466_/Y _11857_/B VGND VGND VPWR VPWR _11813_/B sky130_fd_sc_hd__o22a_1
XFILLER_27_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14525_/X _14529_/X _14525_/X _14529_/X VGND VGND VPWR VPWR _14531_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12791_ _12786_/A _12786_/B _12786_/Y VGND VGND VPWR VPWR _12791_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11780_/B VGND VGND VPWR VPWR _11742_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11576_/Y _11672_/X _11576_/Y _11672_/X VGND VGND VPWR VPWR _11676_/B sky130_fd_sc_hd__a2bb2o_1
X_14461_ _14453_/Y _14459_/X _14460_/Y VGND VGND VPWR VPWR _14461_/X sky130_fd_sc_hd__o21a_1
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16200_ _16103_/X _16199_/X _16103_/X _16199_/X VGND VGND VPWR VPWR _16201_/B sky130_fd_sc_hd__o2bb2a_1
X_14392_ _14317_/X _14390_/X _15597_/B VGND VGND VPWR VPWR _14392_/X sky130_fd_sc_hd__o21a_1
X_13412_ _14908_/A _13415_/B VGND VGND VPWR VPWR _13412_/X sky130_fd_sc_hd__and2_1
X_10624_ _12234_/A _11795_/B VGND VGND VPWR VPWR _12917_/A sky130_fd_sc_hd__or2_1
X_16131_ _16205_/A VGND VGND VPWR VPWR _16189_/A sky130_fd_sc_hd__clkbuf_2
X_13343_ _13275_/X _13342_/Y _13275_/X _13342_/Y VGND VGND VPWR VPWR _13344_/B sky130_fd_sc_hd__a2bb2o_1
X_10555_ _10552_/Y _12697_/A _10451_/X _10554_/Y VGND VGND VPWR VPWR _10555_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16062_ _16062_/A _16053_/X VGND VGND VPWR VPWR _16062_/Y sky130_fd_sc_hd__nor2b_1
X_13274_ _13274_/A _13274_/B VGND VGND VPWR VPWR _13274_/Y sky130_fd_sc_hd__nand2_1
X_10486_ _11773_/A _10392_/B _11773_/A _10392_/B VGND VGND VPWR VPWR _10486_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12225_ _12142_/X _12224_/X _12142_/X _12224_/X VGND VGND VPWR VPWR _12226_/B sky130_fd_sc_hd__a2bb2o_1
X_15013_ _11929_/Y _15003_/X _11929_/Y _15003_/X VGND VGND VPWR VPWR _15040_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12156_ _12206_/A _12154_/X _12155_/X VGND VGND VPWR VPWR _12156_/X sky130_fd_sc_hd__o21a_1
XFILLER_78_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11107_ _11107_/A VGND VGND VPWR VPWR _11107_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12087_ _10980_/A _12086_/A _10980_/Y _12176_/B VGND VGND VPWR VPWR _12089_/B sky130_fd_sc_hd__o22a_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15915_ _15972_/A _15972_/B VGND VGND VPWR VPWR _15915_/X sky130_fd_sc_hd__and2_1
X_11038_ _15075_/A VGND VGND VPWR VPWR _13917_/A sky130_fd_sc_hd__buf_1
XFILLER_49_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15846_ _14201_/A _15845_/X _12628_/X VGND VGND VPWR VPWR _15846_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15777_ _15777_/A _16028_/A VGND VGND VPWR VPWR _15777_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12989_ _14464_/A _12932_/B _12932_/Y VGND VGND VPWR VPWR _12989_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14728_ _14728_/A _14728_/B VGND VGND VPWR VPWR _14728_/X sky130_fd_sc_hd__or2_1
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14659_ _15345_/A _14659_/B VGND VGND VPWR VPWR _14659_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16329_ _16296_/Y _16327_/X _16328_/Y VGND VGND VPWR VPWR _16329_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09703_ _09703_/A VGND VGND VPWR VPWR _09723_/A sky130_fd_sc_hd__inv_2
XFILLER_55_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09634_ _09629_/B _09633_/Y _09629_/B _09633_/Y VGND VGND VPWR VPWR _09635_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09565_ _09563_/Y _09564_/X _09563_/Y _09564_/X VGND VGND VPWR VPWR _09999_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08516_ _08516_/A VGND VGND VPWR VPWR _08516_/Y sky130_fd_sc_hd__clkinvlp_2
X_09496_ _09496_/A _09496_/B VGND VGND VPWR VPWR _09496_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08447_ _08447_/A VGND VGND VPWR VPWR _08447_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08378_ input7/X _08235_/B _08238_/B _08465_/A VGND VGND VPWR VPWR _08378_/X sky130_fd_sc_hd__o22a_2
XFILLER_109_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10340_ _08929_/B _10339_/Y _08928_/A _10277_/Y _10445_/A VGND VGND VPWR VPWR _11718_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10271_ _09297_/A _10230_/B _10231_/A VGND VGND VPWR VPWR _10272_/A sky130_fd_sc_hd__o21ai_1
X_12010_ _12070_/A _12070_/B VGND VGND VPWR VPWR _12010_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13961_ _15420_/A _13961_/B VGND VGND VPWR VPWR _13961_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15700_ _15700_/A _15700_/B VGND VGND VPWR VPWR _15991_/A sky130_fd_sc_hd__or2_1
XFILLER_100_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12912_ _12925_/A _12926_/B VGND VGND VPWR VPWR _12912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13892_ _15418_/A _13959_/B VGND VGND VPWR VPWR _13892_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _14910_/A _15524_/B _15524_/Y VGND VGND VPWR VPWR _15633_/A sky130_fd_sc_hd__o21ai_1
XFILLER_104_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12843_ _12843_/A _12843_/B VGND VGND VPWR VPWR _12843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15562_ _15559_/X _15561_/X _15559_/X _15561_/X VGND VGND VPWR VPWR _15562_/X sky130_fd_sc_hd__a2bb2o_1
X_12774_ _12774_/A _12774_/B VGND VGND VPWR VPWR _12774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15493_ _15484_/X _15492_/X _15484_/X _15492_/X VGND VGND VPWR VPWR _15550_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _15205_/A _14513_/B VGND VGND VPWR VPWR _14513_/X sky130_fd_sc_hd__or2_1
X_11725_ _10282_/A _11724_/Y _10902_/B _10347_/A VGND VGND VPWR VPWR _11736_/B sky130_fd_sc_hd__o22a_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _14466_/A _14466_/B VGND VGND VPWR VPWR _14444_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11656_ _11656_/A VGND VGND VPWR VPWR _13988_/A sky130_fd_sc_hd__buf_1
XFILLER_80_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14375_ _14375_/A _14375_/B VGND VGND VPWR VPWR _15661_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11587_ _13139_/A VGND VGND VPWR VPWR _11656_/A sky130_fd_sc_hd__clkinvlp_2
X_10607_ _10526_/X _10606_/Y _10526_/X _10606_/Y VGND VGND VPWR VPWR _10635_/B sky130_fd_sc_hd__a2bb2o_1
X_16114_ _16114_/A _16114_/B VGND VGND VPWR VPWR _16155_/B sky130_fd_sc_hd__or2_1
X_13326_ _14734_/A _13291_/B _13291_/Y VGND VGND VPWR VPWR _13326_/Y sky130_fd_sc_hd__o21ai_1
X_10538_ _11870_/A VGND VGND VPWR VPWR _13632_/A sky130_fd_sc_hd__buf_1
X_16045_ _16004_/Y _16043_/X _16044_/Y VGND VGND VPWR VPWR _16045_/X sky130_fd_sc_hd__o21a_1
X_13257_ _14424_/A VGND VGND VPWR VPWR _14726_/A sky130_fd_sc_hd__buf_1
XFILLER_89_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12208_ _14014_/A _12208_/B VGND VGND VPWR VPWR _12208_/Y sky130_fd_sc_hd__nand2_1
X_10469_ _09312_/A _10254_/B _10255_/A VGND VGND VPWR VPWR _10470_/A sky130_fd_sc_hd__o21ai_1
XFILLER_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13188_ _13188_/A _13188_/B VGND VGND VPWR VPWR _13188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12139_ _12139_/A _12139_/B VGND VGND VPWR VPWR _12139_/X sky130_fd_sc_hd__or2_1
XFILLER_96_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15829_ _15824_/X _15828_/Y _15824_/X _15828_/Y VGND VGND VPWR VPWR _15829_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09350_ _09350_/A VGND VGND VPWR VPWR _09350_/Y sky130_fd_sc_hd__inv_2
X_08301_ _08400_/B VGND VGND VPWR VPWR _08663_/B sky130_fd_sc_hd__inv_2
X_09281_ _09255_/X _08963_/Y _09255_/X _08963_/Y VGND VGND VPWR VPWR _10250_/A sky130_fd_sc_hd__o2bb2a_1
X_08232_ _08232_/A VGND VGND VPWR VPWR _08233_/A sky130_fd_sc_hd__buf_1
XFILLER_20_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08996_ _08988_/X _08995_/X _08988_/X _08995_/X VGND VGND VPWR VPWR _08997_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09617_ _09508_/X _09616_/X _09508_/X _09616_/X VGND VGND VPWR VPWR _09974_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09548_ _09648_/A _09546_/Y _09648_/B VGND VGND VPWR VPWR _09548_/X sky130_fd_sc_hd__o21ba_1
X_11510_ _13500_/A _11510_/B VGND VGND VPWR VPWR _11510_/X sky130_fd_sc_hd__and2_1
X_09479_ _09448_/Y _09477_/X _09478_/X VGND VGND VPWR VPWR _09520_/S sky130_fd_sc_hd__o21ai_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12490_ _12483_/X _12489_/Y _12483_/X _12489_/Y VGND VGND VPWR VPWR _12490_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11441_ _11256_/X _11440_/Y _11256_/X _11440_/Y VGND VGND VPWR VPWR _12566_/A sky130_fd_sc_hd__a2bb2o_1
X_11372_ _12308_/A _11372_/B VGND VGND VPWR VPWR _11372_/Y sky130_fd_sc_hd__nand2_1
X_14160_ _14145_/X _14159_/Y _14145_/X _14159_/Y VGND VGND VPWR VPWR _14161_/B sky130_fd_sc_hd__a2bb2oi_1
X_13111_ _15255_/A _13111_/B VGND VGND VPWR VPWR _13111_/Y sky130_fd_sc_hd__nand2_1
X_10323_ _11779_/A VGND VGND VPWR VPWR _10324_/A sky130_fd_sc_hd__inv_2
XFILLER_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14091_ _14087_/X _14089_/Y _14222_/B VGND VGND VPWR VPWR _14095_/B sky130_fd_sc_hd__o21ai_1
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13042_ _15234_/A _13125_/B VGND VGND VPWR VPWR _13042_/Y sky130_fd_sc_hd__nor2_1
X_10254_ _10254_/A _10254_/B VGND VGND VPWR VPWR _10255_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10185_ _10468_/A _10167_/B _10167_/Y _10461_/A VGND VGND VPWR VPWR _10564_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14993_ _15781_/B VGND VGND VPWR VPWR _15766_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13944_ _13924_/Y _13942_/X _13943_/Y VGND VGND VPWR VPWR _13944_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13875_ _15110_/A _13974_/B VGND VGND VPWR VPWR _13875_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15614_ _15677_/A _15677_/B VGND VGND VPWR VPWR _15614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12826_ _12826_/A _12839_/B VGND VGND VPWR VPWR _12826_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15545_ _15503_/X _15543_/X _15593_/B VGND VGND VPWR VPWR _15545_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12766_/A _12766_/B VGND VGND VPWR VPWR _12757_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11708_ _11708_/A VGND VGND VPWR VPWR _11709_/A sky130_fd_sc_hd__buf_2
X_15476_ _15467_/A _15467_/B _15467_/Y _15475_/X VGND VGND VPWR VPWR _15476_/X sky130_fd_sc_hd__a2bb2o_1
X_12688_ _10980_/A _12671_/A _10980_/Y _12671_/Y VGND VGND VPWR VPWR _12689_/B sky130_fd_sc_hd__o22a_1
XFILLER_128_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11639_ _12864_/A _11639_/B VGND VGND VPWR VPWR _11639_/X sky130_fd_sc_hd__or2_1
X_14427_ _11788_/X _14413_/X _11788_/X _14413_/X VGND VGND VPWR VPWR _14428_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14358_ _13410_/Y _14357_/Y _13410_/A _14357_/A _14352_/A VGND VGND VPWR VPWR _15948_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13309_ _14067_/A _13309_/B VGND VGND VPWR VPWR _13309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14289_ _14166_/Y _14288_/X _14166_/Y _14288_/X VGND VGND VPWR VPWR _14404_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16028_ _16028_/A _16028_/B VGND VGND VPWR VPWR _16028_/X sky130_fd_sc_hd__or2_1
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08850_ _08852_/A VGND VGND VPWR VPWR _09503_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08781_ _08781_/A VGND VGND VPWR VPWR _08781_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09402_ _09817_/B _09707_/B _09401_/Y VGND VGND VPWR VPWR _09404_/A sky130_fd_sc_hd__a21oi_1
XFILLER_111_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09333_ _09452_/A _10130_/A VGND VGND VPWR VPWR _10044_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09264_ _09242_/X _09263_/X _09242_/X _09263_/X VGND VGND VPWR VPWR _09265_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09195_ _09167_/Y _09194_/Y _09167_/Y _09194_/Y VGND VGND VPWR VPWR _09198_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08979_ _08890_/X _08977_/X _11366_/B VGND VGND VPWR VPWR _08979_/X sky130_fd_sc_hd__o21a_1
X_11990_ _11990_/A VGND VGND VPWR VPWR _12077_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_29_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10941_ _09779_/A _09779_/B _09779_/Y VGND VGND VPWR VPWR _10942_/A sky130_fd_sc_hd__o21ai_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13660_ _13698_/A _13698_/B VGND VGND VPWR VPWR _13729_/A sky130_fd_sc_hd__and2_1
XFILLER_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12611_ _12611_/A VGND VGND VPWR VPWR _12611_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10872_ _10872_/A VGND VGND VPWR VPWR _10872_/Y sky130_fd_sc_hd__inv_2
X_13591_ _13578_/X _13590_/Y _13578_/X _13590_/Y VGND VGND VPWR VPWR _13633_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12542_ _13437_/A _12314_/B _12314_/Y VGND VGND VPWR VPWR _12543_/B sky130_fd_sc_hd__o21a_1
X_15330_ _15329_/A _15329_/B _12045_/Y _15329_/Y VGND VGND VPWR VPWR _15330_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_61_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15261_ _15261_/A _15261_/B VGND VGND VPWR VPWR _15261_/Y sky130_fd_sc_hd__nand2_1
X_12473_ _12471_/Y _12472_/Y _12471_/Y _12472_/Y VGND VGND VPWR VPWR _12473_/X sky130_fd_sc_hd__o2bb2a_1
X_14212_ _14230_/A _14212_/B VGND VGND VPWR VPWR _15872_/A sky130_fd_sc_hd__or2_1
X_11424_ _14083_/A _11424_/B VGND VGND VPWR VPWR _11424_/Y sky130_fd_sc_hd__nor2_1
X_15192_ _15153_/X _15191_/Y _15153_/X _15191_/Y VGND VGND VPWR VPWR _15193_/B sky130_fd_sc_hd__a2bb2o_1
XANTENNA_8 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14143_ _14143_/A VGND VGND VPWR VPWR _14407_/A sky130_fd_sc_hd__inv_2
X_11355_ _14063_/A _11355_/B VGND VGND VPWR VPWR _11355_/Y sky130_fd_sc_hd__nand2_1
X_14074_ _13996_/X _14073_/Y _13996_/X _14073_/Y VGND VGND VPWR VPWR _14074_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11286_ _09995_/A _09664_/B _09664_/Y VGND VGND VPWR VPWR _11286_/X sky130_fd_sc_hd__o21a_1
X_10306_ _10182_/A _10305_/A _10182_/Y _10305_/Y _10462_/A VGND VGND VPWR VPWR _10369_/B
+ sky130_fd_sc_hd__a221o_1
X_13025_ _14411_/A _13025_/B VGND VGND VPWR VPWR _13025_/X sky130_fd_sc_hd__or2_1
XFILLER_4_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ _11577_/A _10237_/B VGND VGND VPWR VPWR _10237_/X sky130_fd_sc_hd__or2_1
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10168_ _10112_/A _10112_/B _10113_/A VGND VGND VPWR VPWR _10251_/A sky130_fd_sc_hd__a21bo_1
X_14976_ _14976_/A _14976_/B VGND VGND VPWR VPWR _14976_/Y sky130_fd_sc_hd__nor2_1
X_10099_ _10099_/A _10099_/B VGND VGND VPWR VPWR _10110_/A sky130_fd_sc_hd__or2_1
X_13927_ _13840_/X _13926_/Y _13840_/X _13926_/Y VGND VGND VPWR VPWR _13941_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13858_ _13802_/Y _13856_/X _13857_/Y VGND VGND VPWR VPWR _13858_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13789_ _15113_/A _13864_/B _13788_/Y VGND VGND VPWR VPWR _13789_/Y sky130_fd_sc_hd__o21ai_1
X_12809_ _12774_/A _12774_/B _12774_/Y VGND VGND VPWR VPWR _12809_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15528_ _15477_/X _15527_/Y _15477_/X _15527_/Y VGND VGND VPWR VPWR _15624_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15459_ _15459_/A _15404_/X VGND VGND VPWR VPWR _15459_/X sky130_fd_sc_hd__or2b_1
XFILLER_128_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09951_ _10216_/A VGND VGND VPWR VPWR _09951_/Y sky130_fd_sc_hd__inv_2
X_08902_ _09551_/A _08596_/A _08598_/A VGND VGND VPWR VPWR _08902_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _09882_/A _09882_/B VGND VGND VPWR VPWR _09883_/B sky130_fd_sc_hd__or2_1
XFILLER_97_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _09228_/A VGND VGND VPWR VPWR _10018_/A sky130_fd_sc_hd__buf_1
XFILLER_111_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _09330_/A _09476_/B _08709_/Y VGND VGND VPWR VPWR _08765_/A sky130_fd_sc_hd__a21oi_2
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08695_ _08871_/A _08693_/X _08871_/B VGND VGND VPWR VPWR _08695_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_26_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09316_ _09262_/A _09262_/B _09262_/X _10801_/A VGND VGND VPWR VPWR _09329_/A sky130_fd_sc_hd__a22o_1
X_09247_ _09247_/A VGND VGND VPWR VPWR _09262_/A sky130_fd_sc_hd__inv_2
X_09178_ _09527_/B _09155_/B _09156_/B VGND VGND VPWR VPWR _09179_/A sky130_fd_sc_hd__a21bo_1
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput34 _16472_/Q VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__clkbuf_2
X_11140_ _12176_/A _11140_/B VGND VGND VPWR VPWR _11140_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11071_ _12137_/A VGND VGND VPWR VPWR _14429_/A sky130_fd_sc_hd__buf_1
XFILLER_88_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10022_ _09251_/A _10125_/A _10065_/B _10021_/X VGND VGND VPWR VPWR _10022_/X sky130_fd_sc_hd__o22a_1
X_14830_ _15351_/A _14830_/B VGND VGND VPWR VPWR _14830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11973_ _11951_/Y _11971_/X _11972_/Y VGND VGND VPWR VPWR _11973_/X sky130_fd_sc_hd__o21a_1
X_14761_ _15181_/A _14761_/B VGND VGND VPWR VPWR _14761_/X sky130_fd_sc_hd__or2_1
XFILLER_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14692_ _14738_/A _14738_/B VGND VGND VPWR VPWR _14780_/A sky130_fd_sc_hd__and2_1
X_10924_ _10924_/A VGND VGND VPWR VPWR _14610_/A sky130_fd_sc_hd__buf_1
X_13712_ _13712_/A _13712_/B VGND VGND VPWR VPWR _13781_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16431_ _16437_/D _16419_/B _16445_/B VGND VGND VPWR VPWR _16431_/Y sky130_fd_sc_hd__o21ai_1
X_10855_ _10921_/A _10922_/B VGND VGND VPWR VPWR _11020_/A sky130_fd_sc_hd__and2_1
X_13643_ _13705_/A VGND VGND VPWR VPWR _15119_/A sky130_fd_sc_hd__buf_1
X_16362_ _16357_/X _16465_/Q _16358_/X _16407_/D _16361_/X VGND VGND VPWR VPWR _16465_/D
+ sky130_fd_sc_hd__o221a_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13574_ _13571_/X _13572_/X _13606_/B VGND VGND VPWR VPWR _13574_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12525_ _12524_/A _12524_/B _12524_/Y _11710_/X VGND VGND VPWR VPWR _12634_/A sky130_fd_sc_hd__o211a_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15313_ _15276_/X _15312_/Y _15276_/X _15312_/Y VGND VGND VPWR VPWR _15339_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ _10784_/Y _10785_/Y _10705_/Y VGND VGND VPWR VPWR _10939_/A sky130_fd_sc_hd__o21ai_1
X_16293_ _16330_/A _16330_/B VGND VGND VPWR VPWR _16293_/Y sky130_fd_sc_hd__nor2_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15244_ _15190_/A _15190_/B _15190_/Y VGND VGND VPWR VPWR _15244_/Y sky130_fd_sc_hd__o21ai_1
X_12456_ _12955_/A _12456_/B VGND VGND VPWR VPWR _12456_/Y sky130_fd_sc_hd__nor2_1
X_15175_ _15556_/A _15556_/B _15174_/Y VGND VGND VPWR VPWR _15175_/Y sky130_fd_sc_hd__o21ai_1
X_12387_ _12437_/B _12386_/Y _12437_/B _12386_/Y VGND VGND VPWR VPWR _12442_/B sky130_fd_sc_hd__o2bb2a_1
X_11407_ _11407_/A VGND VGND VPWR VPWR _11407_/Y sky130_fd_sc_hd__inv_2
X_14126_ _14126_/A VGND VGND VPWR VPWR _14126_/Y sky130_fd_sc_hd__inv_2
X_11338_ _13785_/A _11506_/B _13785_/A _11506_/B VGND VGND VPWR VPWR _11338_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14057_ _14057_/A _14057_/B VGND VGND VPWR VPWR _14057_/X sky130_fd_sc_hd__or2_1
X_11269_ _11177_/A _11095_/X _11176_/X VGND VGND VPWR VPWR _11269_/X sky130_fd_sc_hd__o21a_1
X_13008_ _13008_/A VGND VGND VPWR VPWR _13009_/A sky130_fd_sc_hd__buf_1
XFILLER_79_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14959_ _14831_/X _14958_/Y _14854_/Y VGND VGND VPWR VPWR _14959_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08480_ input26/X input10/X VGND VGND VPWR VPWR _08480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09101_ _09101_/A VGND VGND VPWR VPWR _10102_/B sky130_fd_sc_hd__inv_2
X_09032_ _09547_/B _09032_/B VGND VGND VPWR VPWR _09033_/B sky130_fd_sc_hd__or2_1
XFILLER_132_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09934_ _09863_/X _09932_/X _09863_/X _09932_/X VGND VGND VPWR VPWR _09934_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_131_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09865_ _08904_/X _08597_/A _09455_/Y _09812_/X VGND VGND VPWR VPWR _09865_/X sky130_fd_sc_hd__o22a_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08816_ _10016_/A VGND VGND VPWR VPWR _08819_/A sky130_fd_sc_hd__buf_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09796_ _10621_/A VGND VGND VPWR VPWR _09797_/A sky130_fd_sc_hd__clkbuf_2
X_08747_ _08708_/Y _08745_/Y _08746_/X VGND VGND VPWR VPWR _09340_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08678_ _08678_/A VGND VGND VPWR VPWR _08678_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10602_/Y _10637_/Y _10639_/Y VGND VGND VPWR VPWR _10641_/A sky130_fd_sc_hd__o21ai_1
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10571_ _10571_/A _10571_/B VGND VGND VPWR VPWR _10571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12310_ _12246_/X _12309_/Y _12246_/X _12309_/Y VGND VGND VPWR VPWR _12311_/B sky130_fd_sc_hd__a2bb2o_1
X_13290_ _13290_/A VGND VGND VPWR VPWR _13290_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12241_ _12229_/A _12229_/B _12229_/Y _12240_/X VGND VGND VPWR VPWR _12241_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12172_ _12172_/A VGND VGND VPWR VPWR _12263_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_122_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11123_ _11122_/Y _10947_/X _10994_/Y VGND VGND VPWR VPWR _11123_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15931_ _15894_/A _15894_/B _15894_/Y VGND VGND VPWR VPWR _15931_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11054_ _13925_/A _11080_/B VGND VGND VPWR VPWR _11236_/A sky130_fd_sc_hd__and2_1
XFILLER_49_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10005_ _09963_/A _09962_/Y _09963_/Y _09962_/A _10445_/A VGND VGND VPWR VPWR _11713_/A
+ sky130_fd_sc_hd__o221a_1
X_15862_ _15900_/A _15900_/B VGND VGND VPWR VPWR _15862_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15793_ _15669_/A _15669_/B _15669_/Y VGND VGND VPWR VPWR _15793_/Y sky130_fd_sc_hd__o21ai_1
X_14813_ _14721_/A _14721_/B _14721_/Y VGND VGND VPWR VPWR _14813_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14744_ _14744_/A VGND VGND VPWR VPWR _15351_/A sky130_fd_sc_hd__buf_1
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11956_ _11897_/A _11955_/Y _11897_/A _11955_/Y VGND VGND VPWR VPWR _11968_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10907_ _10907_/A _11413_/A VGND VGND VPWR VPWR _12043_/B sky130_fd_sc_hd__or2_1
XFILLER_60_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16414_ _16437_/D _16473_/Q VGND VGND VPWR VPWR _16415_/A sky130_fd_sc_hd__or2_1
X_11887_ _11837_/X _11886_/Y _11837_/X _11886_/Y VGND VGND VPWR VPWR _11895_/B sky130_fd_sc_hd__a2bb2o_1
X_14675_ _14670_/X _14674_/X _14670_/X _14674_/X VGND VGND VPWR VPWR _14676_/B sky130_fd_sc_hd__a2bb2o_1
X_13626_ _13598_/Y _13623_/Y _13625_/Y VGND VGND VPWR VPWR _13627_/A sky130_fd_sc_hd__o21ai_1
X_10838_ _10799_/X _10837_/X _10799_/X _10837_/X VGND VGND VPWR VPWR _10946_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16345_ _16338_/A _16338_/B _16338_/Y VGND VGND VPWR VPWR _16345_/Y sky130_fd_sc_hd__o21ai_1
X_10769_ _13101_/A _10769_/B VGND VGND VPWR VPWR _10769_/X sky130_fd_sc_hd__or2_1
X_13557_ _15034_/A _13521_/B _13521_/Y VGND VGND VPWR VPWR _13557_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16276_ _16277_/A _16277_/B VGND VGND VPWR VPWR _16276_/X sky130_fd_sc_hd__and2_1
X_12508_ _12508_/A _12508_/B VGND VGND VPWR VPWR _12508_/Y sky130_fd_sc_hd__nand2_1
X_13488_ _10962_/Y _11999_/A _10832_/Y _13487_/X VGND VGND VPWR VPWR _13488_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15227_ _15184_/A _15184_/B _15184_/Y _15226_/X VGND VGND VPWR VPWR _15227_/X sky130_fd_sc_hd__a2bb2o_1
X_12439_ _12439_/A _12439_/B VGND VGND VPWR VPWR _12439_/X sky130_fd_sc_hd__or2_1
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15158_ _15113_/A _15113_/B _15113_/Y _15157_/X VGND VGND VPWR VPWR _15158_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14109_ _15455_/A _14023_/B _14108_/A _14023_/B VGND VGND VPWR VPWR _14109_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15089_ _12139_/A _15084_/B _15084_/Y _15088_/X VGND VGND VPWR VPWR _15089_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09650_ _09975_/A _09650_/B VGND VGND VPWR VPWR _09650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08601_ _08650_/A _08601_/B VGND VGND VPWR VPWR _09456_/B sky130_fd_sc_hd__or2_1
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09581_ _09514_/X _09580_/X _09514_/X _09580_/X VGND VGND VPWR VPWR _09992_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08532_ _08532_/A _08532_/B VGND VGND VPWR VPWR _09861_/A sky130_fd_sc_hd__or2_2
XFILLER_63_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08463_ _08521_/B _08459_/Y _09448_/A VGND VGND VPWR VPWR _08464_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08394_ _08662_/A _08394_/B VGND VGND VPWR VPWR _08395_/A sky130_fd_sc_hd__or2_2
X_09015_ _08778_/A _09014_/Y _08555_/B VGND VGND VPWR VPWR _09015_/X sky130_fd_sc_hd__o21ba_1
XFILLER_132_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09917_ _10949_/B _09917_/B VGND VGND VPWR VPWR _09918_/B sky130_fd_sc_hd__nand2b_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09848_ _09848_/A _09848_/B VGND VGND VPWR VPWR _09848_/X sky130_fd_sc_hd__and2_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09779_ _09779_/A _09779_/B VGND VGND VPWR VPWR _09779_/Y sky130_fd_sc_hd__nand2_1
X_12790_ _12789_/A _12789_/B _12789_/Y VGND VGND VPWR VPWR _12790_/X sky130_fd_sc_hd__a21o_1
X_11810_ _11810_/A VGND VGND VPWR VPWR _11857_/B sky130_fd_sc_hd__inv_2
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11741_ _11745_/B _11740_/Y _11745_/B _11740_/Y VGND VGND VPWR VPWR _11780_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11671_/A _15433_/A _11671_/Y VGND VGND VPWR VPWR _11672_/X sky130_fd_sc_hd__a21o_1
X_14460_ _14460_/A _14460_/B VGND VGND VPWR VPWR _14460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13411_ _14901_/A _13407_/B _13407_/X _13410_/Y VGND VGND VPWR VPWR _13415_/B sky130_fd_sc_hd__o22a_1
X_14391_ _15962_/A _14391_/B VGND VGND VPWR VPWR _15597_/B sky130_fd_sc_hd__or2_1
X_10623_ _10623_/A _10625_/C VGND VGND VPWR VPWR _10626_/A sky130_fd_sc_hd__nor2_1
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16130_ _16243_/A VGND VGND VPWR VPWR _16205_/A sky130_fd_sc_hd__buf_6
X_13342_ _14724_/A _13276_/B _13276_/Y VGND VGND VPWR VPWR _13342_/Y sky130_fd_sc_hd__o21ai_1
X_10554_ _10554_/A _11813_/A VGND VGND VPWR VPWR _10554_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16061_ _16123_/A _16123_/B VGND VGND VPWR VPWR _16061_/X sky130_fd_sc_hd__and2_1
X_13273_ _14721_/A _13272_/B _11415_/X _13272_/Y VGND VGND VPWR VPWR _13273_/X sky130_fd_sc_hd__o2bb2a_1
X_10485_ _11844_/A VGND VGND VPWR VPWR _13624_/A sky130_fd_sc_hd__buf_1
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12224_ _12224_/A _12143_/X VGND VGND VPWR VPWR _12224_/X sky130_fd_sc_hd__or2b_1
X_15012_ _15042_/A _15042_/B VGND VGND VPWR VPWR _15061_/A sky130_fd_sc_hd__and2_1
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12155_ _13897_/A _12155_/B VGND VGND VPWR VPWR _12155_/X sky130_fd_sc_hd__or2_1
XFILLER_69_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11106_ _11106_/A VGND VGND VPWR VPWR _11106_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12086_ _12086_/A VGND VGND VPWR VPWR _12176_/B sky130_fd_sc_hd__inv_2
X_15914_ _15909_/Y _15913_/Y _15909_/Y _15913_/Y VGND VGND VPWR VPWR _15972_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11037_ _12845_/A VGND VGND VPWR VPWR _15075_/A sky130_fd_sc_hd__clkbuf_2
X_15845_ _14207_/A _15844_/X _12626_/X VGND VGND VPWR VPWR _15845_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15776_ _16084_/A VGND VGND VPWR VPWR _15785_/A sky130_fd_sc_hd__inv_2
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12988_ _13692_/A VGND VGND VPWR VPWR _14488_/A sky130_fd_sc_hd__inv_2
X_14727_ _14804_/A _14725_/Y _14726_/X VGND VGND VPWR VPWR _14727_/X sky130_fd_sc_hd__o21a_1
X_11939_ _11980_/A _11980_/B VGND VGND VPWR VPWR _11939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14658_ _14617_/Y _14656_/X _14657_/Y VGND VGND VPWR VPWR _14658_/X sky130_fd_sc_hd__o21a_1
X_13609_ _13609_/A VGND VGND VPWR VPWR _13609_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16328_ _16328_/A _16328_/B VGND VGND VPWR VPWR _16328_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14589_ _15243_/A VGND VGND VPWR VPWR _14664_/A sky130_fd_sc_hd__buf_1
X_16259_ _16202_/Y _16256_/X _16258_/Y VGND VGND VPWR VPWR _16259_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09702_ _09695_/A _09695_/B _09698_/A VGND VGND VPWR VPWR _09970_/A sky130_fd_sc_hd__a21bo_1
XFILLER_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09633_ _08679_/A _09028_/A _09540_/X VGND VGND VPWR VPWR _09633_/Y sky130_fd_sc_hd__o21ai_1
X_09564_ _09478_/A _09518_/B _09478_/A _09518_/B VGND VGND VPWR VPWR _09564_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08515_ _09561_/A _08989_/A _08514_/Y VGND VGND VPWR VPWR _08515_/X sky130_fd_sc_hd__a21o_1
X_09495_ _08814_/X _09465_/X _08814_/X _09465_/X VGND VGND VPWR VPWR _09496_/B sky130_fd_sc_hd__o2bb2a_1
X_08446_ _08446_/A VGND VGND VPWR VPWR _08446_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08377_ _08242_/A input6/X _08307_/B _08460_/A VGND VGND VPWR VPWR _08465_/A sky130_fd_sc_hd__o22a_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10270_ _11745_/A VGND VGND VPWR VPWR _10325_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13960_ _13892_/Y _13958_/X _13959_/Y VGND VGND VPWR VPWR _13960_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12911_ _12838_/X _12910_/Y _12838_/X _12910_/Y VGND VGND VPWR VPWR _12926_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ _15673_/A _15673_/B VGND VGND VPWR VPWR _15630_/Y sky130_fd_sc_hd__nor2_1
X_13891_ _13858_/X _13890_/Y _13858_/X _13890_/Y VGND VGND VPWR VPWR _13959_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12842_ _12823_/Y _12840_/X _12841_/Y VGND VGND VPWR VPWR _12842_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12773_ _12748_/Y _12771_/X _12772_/Y VGND VGND VPWR VPWR _12773_/X sky130_fd_sc_hd__o21a_1
X_15561_ _12428_/A _12429_/B _15560_/Y _15161_/A VGND VGND VPWR VPWR _15561_/X sky130_fd_sc_hd__o22a_1
XFILLER_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15440_/A _15440_/B _15440_/A _15440_/B VGND VGND VPWR VPWR _15492_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14560_/A _14510_/X _14511_/X VGND VGND VPWR VPWR _14512_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11724_ _11724_/A _11724_/B VGND VGND VPWR VPWR _11724_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11656_/A _11657_/B VGND VGND VPWR VPWR _11655_/X sky130_fd_sc_hd__and2_1
X_14443_ _14434_/X _14442_/X _14434_/X _14442_/X VGND VGND VPWR VPWR _14466_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14374_ _14374_/A VGND VGND VPWR VPWR _14374_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10606_ _13605_/A _10527_/B _10527_/Y VGND VGND VPWR VPWR _10606_/Y sky130_fd_sc_hd__o21ai_1
X_11586_ _11586_/A _11586_/B VGND VGND VPWR VPWR _13139_/A sky130_fd_sc_hd__or2_2
XFILLER_127_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16113_ _16070_/X _16111_/X _16163_/B VGND VGND VPWR VPWR _16113_/X sky130_fd_sc_hd__o21a_1
X_13325_ _13364_/A _13364_/B VGND VGND VPWR VPWR _13387_/A sky130_fd_sc_hd__and2_1
X_10537_ _12936_/A VGND VGND VPWR VPWR _11870_/A sky130_fd_sc_hd__inv_2
X_16044_ _16044_/A _16044_/B VGND VGND VPWR VPWR _16044_/Y sky130_fd_sc_hd__nand2_1
X_13256_ _15078_/A VGND VGND VPWR VPWR _14424_/A sky130_fd_sc_hd__inv_2
X_10468_ _10468_/A VGND VGND VPWR VPWR _10468_/Y sky130_fd_sc_hd__inv_2
X_12207_ _12154_/X _12206_/X _12154_/X _12206_/X VGND VGND VPWR VPWR _12208_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_97_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13187_ _13174_/Y _13185_/X _13186_/Y VGND VGND VPWR VPWR _13187_/X sky130_fd_sc_hd__o21a_1
X_10399_ _10359_/X _10398_/X _10359_/X _10398_/X VGND VGND VPWR VPWR _10400_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12138_ _13935_/A _13935_/B _12136_/X _12235_/A VGND VGND VPWR VPWR _12138_/X sky130_fd_sc_hd__a31o_1
XFILLER_97_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12069_ _12068_/Y _11979_/X _12013_/Y VGND VGND VPWR VPWR _12069_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15828_ _15826_/Y _15827_/X _15826_/Y _15827_/X VGND VGND VPWR VPWR _15828_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_65_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15759_ _16101_/A VGND VGND VPWR VPWR _16104_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09280_ _09239_/Y _09279_/X _09239_/Y _09279_/X VGND VGND VPWR VPWR _09946_/A sky130_fd_sc_hd__a2bb2o_2
X_08300_ _08298_/X _08299_/X _08298_/X _08299_/X VGND VGND VPWR VPWR _08400_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08995_ _08990_/Y _08994_/X _08990_/Y _08994_/X VGND VGND VPWR VPWR _08995_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09616_ _09498_/A _09498_/B _09498_/Y VGND VGND VPWR VPWR _09616_/X sky130_fd_sc_hd__a21o_1
X_09547_ _09547_/A _09547_/B VGND VGND VPWR VPWR _09648_/B sky130_fd_sc_hd__and2_1
XFILLER_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09478_ _09478_/A _09478_/B VGND VGND VPWR VPWR _09478_/X sky130_fd_sc_hd__or2_1
XFILLER_12_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08429_ _08429_/A VGND VGND VPWR VPWR _08429_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11440_ _14031_/A _11225_/B _11225_/Y VGND VGND VPWR VPWR _11440_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11371_ _11261_/X _11370_/Y _11261_/X _11370_/Y VGND VGND VPWR VPWR _11372_/B sky130_fd_sc_hd__a2bb2o_1
X_14090_ _14090_/A _14090_/B VGND VGND VPWR VPWR _14222_/B sky130_fd_sc_hd__or2_1
X_13110_ _13082_/Y _13108_/X _13109_/Y VGND VGND VPWR VPWR _13110_/X sky130_fd_sc_hd__o21a_1
X_10322_ _10344_/B _10322_/B VGND VGND VPWR VPWR _11779_/A sky130_fd_sc_hd__or2_2
X_13041_ _13034_/X _13040_/X _13034_/X _13040_/X VGND VGND VPWR VPWR _13125_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10253_ _10250_/Y _10251_/Y _10252_/Y VGND VGND VPWR VPWR _10254_/B sky130_fd_sc_hd__o21ai_2
XFILLER_133_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10184_ _10251_/A _10170_/B _10170_/Y _10377_/A VGND VGND VPWR VPWR _10461_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14992_ _14975_/X _14991_/X _14975_/X _14991_/X VGND VGND VPWR VPWR _15781_/B sky130_fd_sc_hd__a2bb2oi_4
XFILLER_87_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13943_ _15402_/A _13943_/B VGND VGND VPWR VPWR _13943_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13874_ _13868_/X _13873_/X _13868_/X _13873_/X VGND VGND VPWR VPWR _13974_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15613_ _14386_/X _15612_/Y _14386_/X _15612_/Y VGND VGND VPWR VPWR _15677_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12825_ _12763_/Y _12824_/Y _12763_/Y _12824_/Y VGND VGND VPWR VPWR _12839_/B sky130_fd_sc_hd__a2bb2o_1
X_15544_ _15544_/A _15544_/B VGND VGND VPWR VPWR _15593_/B sky130_fd_sc_hd__or2_1
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12710_/X _12755_/X _12710_/X _12755_/X VGND VGND VPWR VPWR _12766_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15475_ _15470_/A _15470_/B _15470_/Y _15474_/X VGND VGND VPWR VPWR _15475_/X sky130_fd_sc_hd__a2bb2o_1
X_11707_ _11680_/X _11706_/X _11680_/X _11706_/X VGND VGND VPWR VPWR _11708_/A sky130_fd_sc_hd__a2bb2oi_4
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _12687_/A _12687_/B VGND VGND VPWR VPWR _12687_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14426_ _15081_/A _14426_/B VGND VGND VPWR VPWR _14426_/X sky130_fd_sc_hd__and2_1
X_11638_ _12864_/A _11639_/B VGND VGND VPWR VPWR _11640_/A sky130_fd_sc_hd__and2_1
XFILLER_128_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14357_ _14357_/A VGND VGND VPWR VPWR _14357_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_116_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11569_ _11569_/A _11569_/B VGND VGND VPWR VPWR _11569_/Y sky130_fd_sc_hd__nand2_1
X_13308_ _13210_/Y _13307_/X _13210_/Y _13307_/X VGND VGND VPWR VPWR _13309_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14288_ _14172_/X _14286_/X _14294_/B VGND VGND VPWR VPWR _14288_/X sky130_fd_sc_hd__o21a_1
X_16027_ _16027_/A _16027_/B VGND VGND VPWR VPWR _16027_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13239_ _13195_/X _13238_/Y _13195_/X _13238_/Y VGND VGND VPWR VPWR _13291_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08780_ _09332_/A _09472_/B _08711_/Y VGND VGND VPWR VPWR _08781_/A sky130_fd_sc_hd__a21oi_2
XFILLER_111_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09401_ _09401_/A _09707_/B VGND VGND VPWR VPWR _09401_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09332_ _09332_/A _09332_/B VGND VGND VPWR VPWR _10041_/A sky130_fd_sc_hd__nor2_1
X_09263_ _09467_/B _09857_/A _09212_/A VGND VGND VPWR VPWR _09263_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09194_ _09340_/A _09161_/Y _09341_/A VGND VGND VPWR VPWR _09194_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08978_ _08978_/A _08978_/B VGND VGND VPWR VPWR _11366_/B sky130_fd_sc_hd__or2_1
X_10940_ _10938_/Y _10939_/Y _10842_/Y VGND VGND VPWR VPWR _11116_/A sky130_fd_sc_hd__o21ai_1
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12610_ _12610_/A VGND VGND VPWR VPWR _12611_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10871_ _09415_/A _09415_/B _09415_/Y VGND VGND VPWR VPWR _10872_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13590_ _13551_/A _13551_/B _13552_/A VGND VGND VPWR VPWR _13590_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12541_ _12540_/A _12540_/B _12540_/Y _11710_/A VGND VGND VPWR VPWR _12630_/A sky130_fd_sc_hd__o211a_1
XFILLER_61_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15260_ _15219_/X _15259_/Y _15219_/X _15259_/Y VGND VGND VPWR VPWR _15261_/B sky130_fd_sc_hd__a2bb2o_1
X_12472_ _13972_/A _12449_/B _12449_/Y _12452_/X VGND VGND VPWR VPWR _12472_/Y sky130_fd_sc_hd__o2bb2ai_1
X_11423_ _13405_/A _13405_/B _12607_/B _11422_/X VGND VGND VPWR VPWR _11424_/B sky130_fd_sc_hd__a31o_1
X_14211_ _14099_/Y _14210_/X _14099_/Y _14210_/X VGND VGND VPWR VPWR _14212_/B sky130_fd_sc_hd__a2bb2oi_1
X_15191_ _15125_/A _15125_/B _15125_/Y VGND VGND VPWR VPWR _15191_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_9 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ _14143_/A _14144_/A VGND VGND VPWR VPWR _14142_/Y sky130_fd_sc_hd__nor2_1
X_11354_ _11269_/X _11353_/X _11269_/X _11353_/X VGND VGND VPWR VPWR _11355_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14073_ _13998_/X _14072_/X _13998_/X _14072_/X VGND VGND VPWR VPWR _14073_/Y sky130_fd_sc_hd__a2bb2oi_1
X_11285_ _12195_/A _11170_/B _11170_/Y _11110_/X VGND VGND VPWR VPWR _11285_/X sky130_fd_sc_hd__a2bb2o_1
X_10305_ _10305_/A VGND VGND VPWR VPWR _10305_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13024_ _13070_/A _13022_/X _13023_/X VGND VGND VPWR VPWR _13024_/X sky130_fd_sc_hd__o21a_1
X_10236_ _10234_/Y _10235_/X _10175_/Y VGND VGND VPWR VPWR _10236_/Y sky130_fd_sc_hd__o21ai_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10167_ _10167_/A _10167_/B VGND VGND VPWR VPWR _10167_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14975_ _14970_/Y _14974_/X _14970_/Y _14974_/X VGND VGND VPWR VPWR _14975_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10098_ _10098_/A _10098_/B VGND VGND VPWR VPWR _10099_/A sky130_fd_sc_hd__or2_1
X_13926_ _14634_/A _13841_/B _13841_/Y VGND VGND VPWR VPWR _13926_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13857_ _14663_/A _13857_/B VGND VGND VPWR VPWR _13857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13788_ _13788_/A _13864_/B VGND VGND VPWR VPWR _13788_/Y sky130_fd_sc_hd__nand2_1
X_12808_ _12851_/A _12851_/B VGND VGND VPWR VPWR _12808_/Y sky130_fd_sc_hd__nor2_1
X_15527_ _15461_/A _15461_/B _15461_/Y VGND VGND VPWR VPWR _15527_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _12778_/A _12778_/B VGND VGND VPWR VPWR _12739_/Y sky130_fd_sc_hd__nor2_1
X_15458_ _15458_/A _15458_/B VGND VGND VPWR VPWR _15458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14409_ _14409_/A VGND VGND VPWR VPWR _15347_/A sky130_fd_sc_hd__buf_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15389_ _15400_/A _15400_/B VGND VGND VPWR VPWR _15465_/A sky130_fd_sc_hd__and2_1
XFILLER_7_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09950_ _11773_/A VGND VGND VPWR VPWR _13559_/A sky130_fd_sc_hd__buf_1
X_08901_ _08974_/A _08974_/B VGND VGND VPWR VPWR _08901_/X sky130_fd_sc_hd__and2_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09865_/X _08806_/Y _09865_/X _08806_/Y VGND VGND VPWR VPWR _09882_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _08831_/X _08725_/Y _08831_/A _08725_/Y VGND VGND VPWR VPWR _08834_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _09331_/A VGND VGND VPWR VPWR _09484_/A sky130_fd_sc_hd__buf_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08694_ _08694_/A _10120_/B VGND VGND VPWR VPWR _08871_/B sky130_fd_sc_hd__and2_1
XFILLER_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09315_ _09268_/A _09268_/B _09268_/X _10664_/A VGND VGND VPWR VPWR _10801_/A sky130_fd_sc_hd__a22o_1
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09246_ _09243_/X _09245_/X _09243_/X _09245_/X VGND VGND VPWR VPWR _09247_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09177_ _09431_/A _09180_/B VGND VGND VPWR VPWR _09177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11070_ _12915_/A VGND VGND VPWR VPWR _12137_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10021_ _09458_/A _10124_/A _10061_/B _10020_/X VGND VGND VPWR VPWR _10021_/X sky130_fd_sc_hd__o22a_1
XFILLER_130_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14760_ _15181_/A _14761_/B VGND VGND VPWR VPWR _14762_/A sky130_fd_sc_hd__and2_1
XFILLER_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11972_ _11972_/A _11972_/B VGND VGND VPWR VPWR _11972_/Y sky130_fd_sc_hd__nand2_1
X_13711_ _13539_/X _13710_/Y _13539_/X _13710_/Y VGND VGND VPWR VPWR _13712_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10923_ _11020_/A _10920_/X _10922_/X VGND VGND VPWR VPWR _10923_/X sky130_fd_sc_hd__o21a_1
X_14691_ _14660_/X _14690_/Y _14660_/X _14690_/Y VGND VGND VPWR VPWR _14738_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16430_ _16416_/Y _16447_/B _16428_/Y _16415_/X _16429_/X VGND VGND VPWR VPWR _16445_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10854_ _10778_/X _10853_/Y _10778_/X _10853_/Y VGND VGND VPWR VPWR _10922_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_72_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13642_ _13586_/Y _13639_/Y _13641_/Y VGND VGND VPWR VPWR _13704_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16361_ _16361_/A VGND VGND VPWR VPWR _16361_/X sky130_fd_sc_hd__buf_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _14428_/A _13573_/B VGND VGND VPWR VPWR _13606_/B sky130_fd_sc_hd__or2_1
X_12524_ _12524_/A _12524_/B VGND VGND VPWR VPWR _12524_/Y sky130_fd_sc_hd__nand2_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ _14581_/A _15255_/B _15255_/Y VGND VGND VPWR VPWR _15312_/Y sky130_fd_sc_hd__o21ai_1
X_10785_ _10785_/A VGND VGND VPWR VPWR _10785_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16292_ _16263_/X _16291_/Y _16263_/X _16291_/Y VGND VGND VPWR VPWR _16330_/B sky130_fd_sc_hd__o2bb2a_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15243_ _15243_/A _15243_/B VGND VGND VPWR VPWR _15243_/Y sky130_fd_sc_hd__nand2_1
X_12455_ _13978_/A _12454_/B _12454_/Y VGND VGND VPWR VPWR _12455_/X sky130_fd_sc_hd__a21o_1
X_11406_ _12331_/A VGND VGND VPWR VPWR _15519_/A sky130_fd_sc_hd__buf_1
X_15174_ _15556_/A _15556_/B VGND VGND VPWR VPWR _15174_/Y sky130_fd_sc_hd__nand2_1
X_12386_ _12786_/A _12385_/B _12385_/Y VGND VGND VPWR VPWR _12386_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14125_ _14125_/A VGND VGND VPWR VPWR _14872_/A sky130_fd_sc_hd__inv_2
X_11337_ _11307_/X _11336_/X _11307_/X _11336_/X VGND VGND VPWR VPWR _11506_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14056_ _14076_/A _14054_/X _14055_/X VGND VGND VPWR VPWR _14056_/X sky130_fd_sc_hd__o21a_1
X_11268_ _14008_/A VGND VGND VPWR VPWR _14063_/A sky130_fd_sc_hd__buf_1
XFILLER_97_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ _12921_/X _13006_/X _12921_/X _13006_/X VGND VGND VPWR VPWR _13010_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10219_ _10454_/A _11232_/A VGND VGND VPWR VPWR _11748_/A sky130_fd_sc_hd__or2_1
X_11199_ _11199_/A VGND VGND VPWR VPWR _11199_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14958_ _15353_/A _14958_/B VGND VGND VPWR VPWR _14958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14889_ _15534_/A _14914_/B VGND VGND VPWR VPWR _14889_/Y sky130_fd_sc_hd__nor2_1
X_13909_ _13909_/A VGND VGND VPWR VPWR _15408_/A sky130_fd_sc_hd__buf_1
XFILLER_63_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09100_ _09709_/A VGND VGND VPWR VPWR _09407_/A sky130_fd_sc_hd__buf_1
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09031_ _09538_/B _09031_/B VGND VGND VPWR VPWR _09032_/B sky130_fd_sc_hd__or2_1
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09933_ _09932_/A _09932_/B _09932_/X VGND VGND VPWR VPWR _09933_/X sky130_fd_sc_hd__a21bo_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09864_ _09863_/A _09863_/B _09863_/X VGND VGND VPWR VPWR _09864_/X sky130_fd_sc_hd__a21bo_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08815_ _08814_/X _08727_/X _08814_/A _08727_/X VGND VGND VPWR VPWR _08817_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09795_ _09196_/Y _09794_/A _09198_/X _09794_/Y VGND VGND VPWR VPWR _10621_/A sky130_fd_sc_hd__o22a_4
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08746_ _10008_/A _09448_/B VGND VGND VPWR VPWR _08746_/X sky130_fd_sc_hd__or2_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08677_ _09234_/A _08677_/B VGND VGND VPWR VPWR _08678_/A sky130_fd_sc_hd__or2_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10570_ _09274_/B _10244_/B _10244_/X VGND VGND VPWR VPWR _10571_/B sky130_fd_sc_hd__a21boi_1
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09229_ _09800_/A VGND VGND VPWR VPWR _09687_/A sky130_fd_sc_hd__inv_2
X_12240_ _13348_/A _12232_/B _12232_/Y _12239_/X VGND VGND VPWR VPWR _12240_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12171_ _12169_/A _12169_/B _12169_/X _12170_/Y VGND VGND VPWR VPWR _12263_/B sky130_fd_sc_hd__a22o_1
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11122_ _12097_/A _11122_/B VGND VGND VPWR VPWR _11122_/Y sky130_fd_sc_hd__nor2_1
X_15930_ _15958_/A _15958_/B VGND VGND VPWR VPWR _15930_/X sky130_fd_sc_hd__and2_1
X_11053_ _10913_/X _11052_/X _10913_/X _11052_/X VGND VGND VPWR VPWR _11080_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15861_ _14189_/X _15847_/X _14189_/X _15847_/X VGND VGND VPWR VPWR _15900_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10004_ _10344_/B VGND VGND VPWR VPWR _10445_/A sky130_fd_sc_hd__inv_2
XFILLER_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14812_ _14812_/A _14812_/B VGND VGND VPWR VPWR _14812_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15792_ _16094_/A _15795_/B VGND VGND VPWR VPWR _15792_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14743_ _14662_/X _14742_/Y _14686_/Y VGND VGND VPWR VPWR _14743_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11955_ _12997_/A _11898_/B _11898_/Y VGND VGND VPWR VPWR _11955_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14674_ _14673_/A _14673_/B _14673_/Y VGND VGND VPWR VPWR _14674_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10906_ _10906_/A VGND VGND VPWR VPWR _11413_/A sky130_fd_sc_hd__clkbuf_2
X_16413_ _16474_/Q VGND VGND VPWR VPWR _16437_/D sky130_fd_sc_hd__inv_2
X_11886_ _11838_/A _11838_/B _11838_/Y VGND VGND VPWR VPWR _11886_/Y sky130_fd_sc_hd__o21ai_1
X_13625_ _15134_/A _13625_/B VGND VGND VPWR VPWR _13625_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10837_ _11009_/A _10953_/B _11009_/A _10953_/B VGND VGND VPWR VPWR _10837_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16344_ _08230_/X _16470_/Q _08233_/X _16392_/A _16343_/X VGND VGND VPWR VPWR _16470_/D
+ sky130_fd_sc_hd__o221a_2
X_10768_ _10768_/A VGND VGND VPWR VPWR _13101_/A sky130_fd_sc_hd__buf_1
X_13556_ _13556_/A VGND VGND VPWR VPWR _13556_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16275_ _16137_/Y _16274_/Y _16137_/Y _16274_/Y VGND VGND VPWR VPWR _16277_/B sky130_fd_sc_hd__a2bb2o_1
X_12507_ _13445_/A _11358_/B _11358_/Y VGND VGND VPWR VPWR _12508_/B sky130_fd_sc_hd__o21a_1
X_13487_ _10810_/Y _11928_/A _10695_/Y _13486_/X VGND VGND VPWR VPWR _13487_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15226_ _15187_/A _15187_/B _15187_/Y _15225_/X VGND VGND VPWR VPWR _15226_/X sky130_fd_sc_hd__a2bb2o_1
X_12438_ _12437_/A _12437_/B _12437_/Y _12385_/B VGND VGND VPWR VPWR _12439_/B sky130_fd_sc_hd__a2bb2o_1
X_10699_ _10668_/X _10698_/X _10668_/X _10698_/X VGND VGND VPWR VPWR _10798_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15157_ _15116_/A _15116_/B _15116_/Y _15156_/X VGND VGND VPWR VPWR _15157_/X sky130_fd_sc_hd__a2bb2o_1
X_12369_ _13785_/A _12369_/B VGND VGND VPWR VPWR _12369_/X sky130_fd_sc_hd__and2_1
XFILLER_4_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14108_ _14108_/A VGND VGND VPWR VPWR _15455_/A sky130_fd_sc_hd__buf_1
X_15088_ _12836_/X _15144_/A _15087_/X VGND VGND VPWR VPWR _15088_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14039_ _14042_/A VGND VGND VPWR VPWR _14812_/A sky130_fd_sc_hd__buf_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08600_ _08599_/A _08348_/Y _08599_/Y _08348_/A VGND VGND VPWR VPWR _08601_/B sky130_fd_sc_hd__o22a_1
XFILLER_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09580_ _09486_/A _09486_/B _09486_/Y VGND VGND VPWR VPWR _09580_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08531_ _09474_/B VGND VGND VPWR VPWR _08692_/A sky130_fd_sc_hd__buf_1
XFILLER_50_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08462_ _08697_/A VGND VGND VPWR VPWR _09448_/A sky130_fd_sc_hd__inv_2
XFILLER_23_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08393_ _08358_/A input18/X _08392_/A _08399_/A _08392_/Y VGND VGND VPWR VPWR _08394_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09014_ _09488_/A _09020_/S _08565_/B VGND VGND VPWR VPWR _09014_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09916_ _10949_/A _10948_/A VGND VGND VPWR VPWR _09917_/B sky130_fd_sc_hd__or2_1
XFILLER_113_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09847_ _10490_/A _09847_/B VGND VGND VPWR VPWR _09848_/B sky130_fd_sc_hd__nand2b_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09778_ _09779_/A _09779_/B VGND VGND VPWR VPWR _09778_/Y sky130_fd_sc_hd__nor2_1
X_08729_ _08729_/A VGND VGND VPWR VPWR _08729_/Y sky130_fd_sc_hd__inv_2
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _10325_/B _11746_/A _11739_/Y VGND VGND VPWR VPWR _11740_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11671_/A _15433_/A VGND VGND VPWR VPWR _11671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13410_ _13410_/A VGND VGND VPWR VPWR _13410_/Y sky130_fd_sc_hd__inv_4
X_14390_ _14323_/X _14388_/X _15605_/B VGND VGND VPWR VPWR _14390_/X sky130_fd_sc_hd__o21a_1
X_10622_ _15212_/A VGND VGND VPWR VPWR _11889_/A sky130_fd_sc_hd__inv_2
X_13341_ _13344_/A VGND VGND VPWR VPWR _15467_/A sky130_fd_sc_hd__buf_1
X_10553_ _11855_/A VGND VGND VPWR VPWR _11813_/A sky130_fd_sc_hd__inv_2
X_16060_ _16054_/X _16059_/Y _16054_/X _16059_/Y VGND VGND VPWR VPWR _16123_/B sky130_fd_sc_hd__a2bb2o_1
X_13272_ _15087_/A _13272_/B VGND VGND VPWR VPWR _13272_/Y sky130_fd_sc_hd__nor2_1
X_10484_ _12932_/A VGND VGND VPWR VPWR _11844_/A sky130_fd_sc_hd__inv_2
X_15011_ _12000_/Y _15004_/X _12000_/Y _15004_/X VGND VGND VPWR VPWR _15042_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12223_ _14028_/A _12223_/B VGND VGND VPWR VPWR _12223_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12154_ _12209_/A _12152_/X _12153_/X VGND VGND VPWR VPWR _12154_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11105_ _09782_/A _09379_/A _09432_/X VGND VGND VPWR VPWR _11106_/A sky130_fd_sc_hd__o21ai_1
X_12085_ _10819_/A _11996_/A _10966_/B _12084_/Y VGND VGND VPWR VPWR _12086_/A sky130_fd_sc_hd__o22a_1
X_15913_ _15978_/A _15978_/B _15912_/Y VGND VGND VPWR VPWR _15913_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11036_ _13559_/A VGND VGND VPWR VPWR _12845_/A sky130_fd_sc_hd__buf_1
XFILLER_134_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15844_ _14213_/A _15843_/X _12624_/X VGND VGND VPWR VPWR _15844_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15775_ _15781_/B _15775_/B VGND VGND VPWR VPWR _16084_/A sky130_fd_sc_hd__or2_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14726_ _14726_/A _14726_/B VGND VGND VPWR VPWR _14726_/X sky130_fd_sc_hd__or2_1
XFILLER_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12987_ _14484_/A _13021_/B VGND VGND VPWR VPWR _13075_/A sky130_fd_sc_hd__and2_1
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11938_ _11913_/X _11937_/Y _11913_/X _11937_/Y VGND VGND VPWR VPWR _11980_/B sky130_fd_sc_hd__a2bb2o_1
X_14657_ _15343_/A _14657_/B VGND VGND VPWR VPWR _14657_/Y sky130_fd_sc_hd__nand2_1
X_11869_ _11849_/X _11868_/X _11849_/X _11868_/X VGND VGND VPWR VPWR _11912_/B sky130_fd_sc_hd__a2bb2o_1
X_14588_ _14538_/Y _14586_/X _14587_/Y VGND VGND VPWR VPWR _14588_/X sky130_fd_sc_hd__o21a_1
X_13608_ _13608_/A _13608_/B VGND VGND VPWR VPWR _13608_/X sky130_fd_sc_hd__and2_1
X_16327_ _16299_/Y _16325_/X _16326_/Y VGND VGND VPWR VPWR _16327_/X sky130_fd_sc_hd__o21a_1
X_13539_ _15044_/A _13506_/B _13506_/Y _13538_/X VGND VGND VPWR VPWR _13539_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16258_ _16324_/A _16258_/B VGND VGND VPWR VPWR _16258_/Y sky130_fd_sc_hd__nand2_1
X_16189_ _16189_/A _16189_/B VGND VGND VPWR VPWR _16260_/A sky130_fd_sc_hd__or2_1
X_15209_ _15143_/A _15143_/B _15143_/Y VGND VGND VPWR VPWR _15209_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09701_ _09701_/A VGND VGND VPWR VPWR _09770_/A sky130_fd_sc_hd__inv_2
XFILLER_110_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09632_ _09632_/A VGND VGND VPWR VPWR _09632_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09563_ _09563_/A VGND VGND VPWR VPWR _09563_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08514_ _09561_/A _08989_/A VGND VGND VPWR VPWR _08514_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09494_ _09494_/A _09494_/B VGND VGND VPWR VPWR _09494_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08445_ _08555_/B _08439_/Y _09332_/A VGND VGND VPWR VPWR _08446_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08376_ input5/X _08245_/B _08312_/B _08375_/X VGND VGND VPWR VPWR _08460_/A sky130_fd_sc_hd__o22a_1
XFILLER_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13890_ _14744_/A _13859_/B _13859_/Y VGND VGND VPWR VPWR _13890_/Y sky130_fd_sc_hd__o21ai_1
X_12910_ _15084_/A _12839_/B _12839_/Y VGND VGND VPWR VPWR _12910_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12841_ _12841_/A _12841_/B VGND VGND VPWR VPWR _12841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12772_ _12772_/A _12772_/B VGND VGND VPWR VPWR _12772_/Y sky130_fd_sc_hd__nand2_1
X_15560_ _15560_/A VGND VGND VPWR VPWR _15560_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15491_ _15552_/A _15552_/B VGND VGND VPWR VPWR _15491_/X sky130_fd_sc_hd__and2_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _15208_/A _14511_/B VGND VGND VPWR VPWR _14511_/X sky130_fd_sc_hd__or2_1
X_11723_ _11723_/A _11723_/B VGND VGND VPWR VPWR _11734_/B sky130_fd_sc_hd__or2_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11654_ _11651_/Y _11653_/X _11651_/Y _11653_/X VGND VGND VPWR VPWR _11657_/B sky130_fd_sc_hd__a2bb2o_1
X_14442_ _14420_/A _14420_/B _14420_/Y VGND VGND VPWR VPWR _14442_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10605_ _09951_/Y _10604_/Y _10216_/X _10604_/A _09797_/A VGND VGND VPWR VPWR _11885_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_128_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14373_ _14247_/A _14370_/X _14372_/Y _14248_/B _14372_/A VGND VGND VPWR VPWR _14374_/A
+ sky130_fd_sc_hd__a32o_1
X_16112_ _16112_/A _16112_/B VGND VGND VPWR VPWR _16163_/B sky130_fd_sc_hd__or2_1
X_11585_ _09440_/X _11584_/X _09440_/X _11584_/X VGND VGND VPWR VPWR _11586_/B sky130_fd_sc_hd__a2bb2o_1
X_13324_ _13293_/A _13323_/Y _13293_/A _13323_/Y VGND VGND VPWR VPWR _13364_/B sky130_fd_sc_hd__a2bb2o_1
X_10536_ _09899_/Y _10535_/X _09898_/X _09901_/B _10794_/A VGND VGND VPWR VPWR _12936_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_10_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16043_ _16007_/Y _16041_/X _16042_/Y VGND VGND VPWR VPWR _16043_/X sky130_fd_sc_hd__o21a_1
X_13255_ _14728_/A _13282_/B VGND VGND VPWR VPWR _13255_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10467_ _10453_/X _10466_/Y _10453_/X _10466_/Y VGND VGND VPWR VPWR _10554_/A sky130_fd_sc_hd__o2bb2a_1
X_12206_ _12206_/A _12155_/X VGND VGND VPWR VPWR _12206_/X sky130_fd_sc_hd__or2b_1
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13186_ _13824_/A _13186_/B VGND VGND VPWR VPWR _13186_/Y sky130_fd_sc_hd__nand2_1
X_10398_ _13524_/A _10319_/B _11713_/A _10319_/B VGND VGND VPWR VPWR _10398_/X sky130_fd_sc_hd__a2bb2o_1
X_12137_ _12137_/A _12137_/B VGND VGND VPWR VPWR _12235_/A sky130_fd_sc_hd__and2_1
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12068_ _12068_/A _12068_/B VGND VGND VPWR VPWR _12068_/Y sky130_fd_sc_hd__nor2_1
X_11019_ _15066_/A VGND VGND VPWR VPWR _13905_/A sky130_fd_sc_hd__buf_1
XFILLER_77_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15827_ _14164_/X _14288_/X _14166_/B VGND VGND VPWR VPWR _15827_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15758_ _15766_/A _15758_/B VGND VGND VPWR VPWR _16101_/A sky130_fd_sc_hd__or2_1
XFILLER_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15689_ _15694_/A _15694_/B VGND VGND VPWR VPWR _15689_/Y sky130_fd_sc_hd__nor2_1
X_14709_ _14648_/X _14708_/Y _14648_/X _14708_/Y VGND VGND VPWR VPWR _14726_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08230_ _08230_/A VGND VGND VPWR VPWR _08230_/X sky130_fd_sc_hd__buf_1
XFILLER_33_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08994_ _08992_/X _08993_/Y _08992_/X _08993_/Y VGND VGND VPWR VPWR _08994_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09615_ _09978_/A _09652_/B VGND VGND VPWR VPWR _09615_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09546_ _09546_/A VGND VGND VPWR VPWR _09546_/Y sky130_fd_sc_hd__inv_2
X_09477_ _09449_/Y _09475_/X _09476_/X VGND VGND VPWR VPWR _09477_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08428_ _09213_/B _08423_/X _08794_/A VGND VGND VPWR VPWR _08428_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08359_ input9/X _08278_/A _08399_/A VGND VGND VPWR VPWR _08359_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11370_ _14059_/A _11188_/B _11188_/Y VGND VGND VPWR VPWR _11370_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10321_ _10216_/X _10320_/Y _10216_/X _10320_/Y VGND VGND VPWR VPWR _10322_/B sky130_fd_sc_hd__o2bb2a_1
X_13040_ _13040_/A _13035_/X VGND VGND VPWR VPWR _13040_/X sky130_fd_sc_hd__or2b_1
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10252_ _10252_/A _10252_/B VGND VGND VPWR VPWR _10252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10183_ _10173_/A _10173_/B _10173_/Y _10182_/Y VGND VGND VPWR VPWR _10377_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_94_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14991_ _14988_/X _14990_/Y _14988_/X _14990_/Y VGND VGND VPWR VPWR _14991_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_78_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13942_ _13928_/Y _13940_/Y _13941_/Y VGND VGND VPWR VPWR _13942_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13873_ _13873_/A _13873_/B VGND VGND VPWR VPWR _13873_/X sky130_fd_sc_hd__or2_1
X_15612_ _14329_/X _15612_/B VGND VGND VPWR VPWR _15612_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_62_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12824_ _12764_/A _12764_/B _12764_/Y VGND VGND VPWR VPWR _12824_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15543_ _15600_/A _15602_/A _15542_/X VGND VGND VPWR VPWR _15543_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12755_ _12704_/A _12704_/B _12704_/A _12704_/B VGND VGND VPWR VPWR _12755_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11706_ _11691_/Y _11705_/Y _11691_/Y _11705_/Y VGND VGND VPWR VPWR _11706_/X sky130_fd_sc_hd__a2bb2o_2
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _15473_/A _15473_/B _12237_/X _15473_/Y VGND VGND VPWR VPWR _15474_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _11152_/A _12673_/A _11152_/Y _12673_/Y VGND VGND VPWR VPWR _12687_/B sky130_fd_sc_hd__o22a_1
X_14425_ _11781_/Y _14415_/A _11781_/Y _14415_/A VGND VGND VPWR VPWR _14426_/B sky130_fd_sc_hd__o2bb2a_1
X_11637_ _11633_/X _11636_/X _11633_/X _11636_/X VGND VGND VPWR VPWR _11639_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14356_ _14906_/A _13407_/B _13407_/X VGND VGND VPWR VPWR _14357_/A sky130_fd_sc_hd__o21ba_1
X_11568_ _13447_/A _11567_/B _11567_/Y VGND VGND VPWR VPWR _11569_/B sky130_fd_sc_hd__o21a_1
X_13307_ _13215_/Y _13305_/Y _13306_/Y VGND VGND VPWR VPWR _13307_/X sky130_fd_sc_hd__o21a_1
X_10519_ _10428_/X _10518_/X _10625_/A _10518_/X VGND VGND VPWR VPWR _10523_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16026_ _14370_/X _15665_/B _14370_/X _15665_/B VGND VGND VPWR VPWR _16027_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14287_ _15910_/A _14287_/B VGND VGND VPWR VPWR _14294_/B sky130_fd_sc_hd__or2_1
X_11499_ _12393_/A VGND VGND VPWR VPWR _12955_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13238_ _13196_/A _13196_/B _13196_/Y VGND VGND VPWR VPWR _13238_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13169_ _15261_/A _13107_/B _13107_/Y VGND VGND VPWR VPWR _13169_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09400_ _09400_/A VGND VGND VPWR VPWR _09707_/B sky130_fd_sc_hd__clkbuf_2
X_09331_ _09331_/A _09331_/B VGND VGND VPWR VPWR _10038_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09262_ _09262_/A _09262_/B VGND VGND VPWR VPWR _09262_/X sky130_fd_sc_hd__or2_1
X_09193_ _09193_/A VGND VGND VPWR VPWR _09193_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08977_ _08896_/X _08975_/X _11373_/B VGND VGND VPWR VPWR _08977_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10870_ _10870_/A _10870_/B VGND VGND VPWR VPWR _10870_/X sky130_fd_sc_hd__and2_1
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09529_ _09529_/A _09529_/B VGND VGND VPWR VPWR _09530_/A sky130_fd_sc_hd__or2_1
XFILLER_101_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12540_ _12540_/A _12540_/B VGND VGND VPWR VPWR _12540_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12471_ _12463_/Y _12470_/X _12463_/Y _12470_/X VGND VGND VPWR VPWR _12471_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_8_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11422_ _13404_/A _11422_/B VGND VGND VPWR VPWR _11422_/X sky130_fd_sc_hd__and2_1
X_14210_ _14100_/A _14100_/B _14100_/Y VGND VGND VPWR VPWR _14210_/X sky130_fd_sc_hd__o21a_1
X_15190_ _15190_/A _15190_/B VGND VGND VPWR VPWR _15190_/Y sky130_fd_sc_hd__nand2_1
X_14141_ _14064_/X _14140_/X _14064_/X _14140_/X VGND VGND VPWR VPWR _14144_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11353_ _11353_/A _11352_/X VGND VGND VPWR VPWR _11353_/X sky130_fd_sc_hd__or2b_1
XFILLER_125_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11284_ _12292_/A VGND VGND VPWR VPWR _11482_/A sky130_fd_sc_hd__inv_2
X_14072_ _13999_/Y _14071_/X _13999_/Y _14071_/X VGND VGND VPWR VPWR _14072_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10304_ _10304_/A1 _10173_/B _10173_/Y VGND VGND VPWR VPWR _10305_/A sky130_fd_sc_hd__a21oi_1
XFILLER_133_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13023_ _14480_/A _13023_/B VGND VGND VPWR VPWR _13023_/X sky130_fd_sc_hd__or2_1
X_10235_ _10235_/A _10235_/B VGND VGND VPWR VPWR _10235_/X sky130_fd_sc_hd__and2_1
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10166_ _10126_/A _10126_/B _10127_/B VGND VGND VPWR VPWR _10167_/B sky130_fd_sc_hd__a21bo_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14974_ _14972_/X _14973_/Y _14972_/X _14973_/Y VGND VGND VPWR VPWR _14974_/X sky130_fd_sc_hd__o2bb2a_1
X_10097_ _11736_/A VGND VGND VPWR VPWR _10213_/A sky130_fd_sc_hd__inv_4
X_13925_ _13925_/A VGND VGND VPWR VPWR _15400_/A sky130_fd_sc_hd__buf_1
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13856_ _13805_/Y _13854_/X _13855_/Y VGND VGND VPWR VPWR _13856_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12807_ _12775_/X _12806_/Y _12775_/X _12806_/Y VGND VGND VPWR VPWR _12851_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10999_ _11116_/A _10998_/Y _11116_/A _10998_/Y VGND VGND VPWR VPWR _11000_/B sky130_fd_sc_hd__a2bb2o_1
X_13787_ _13782_/X _13786_/Y _13782_/X _13786_/Y VGND VGND VPWR VPWR _13864_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15526_ _15529_/A _15529_/B VGND VGND VPWR VPWR _15526_/Y sky130_fd_sc_hd__nor2_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12716_/X _12737_/X _12716_/X _12737_/X VGND VGND VPWR VPWR _12778_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15457_ _15405_/X _15456_/X _15405_/X _15456_/X VGND VGND VPWR VPWR _15458_/B sky130_fd_sc_hd__a2bb2o_1
X_12669_ _12669_/A VGND VGND VPWR VPWR _12669_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14408_ _15440_/A VGND VGND VPWR VPWR _14774_/A sky130_fd_sc_hd__buf_1
XFILLER_30_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15388_ _15332_/X _15387_/X _15332_/X _15387_/X VGND VGND VPWR VPWR _15400_/B sky130_fd_sc_hd__a2bb2o_1
X_14339_ _13424_/Y _14338_/X _13424_/Y _14338_/X VGND VGND VPWR VPWR _14340_/B sky130_fd_sc_hd__a2bb2oi_1
X_16009_ _15957_/X _16008_/Y _15957_/X _16008_/Y VGND VGND VPWR VPWR _16040_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09866_/X _08797_/A _09866_/X _08797_/A VGND VGND VPWR VPWR _09883_/A sky130_fd_sc_hd__a2bb2o_1
X_08900_ _08899_/Y _08862_/X _08899_/Y _08862_/X VGND VGND VPWR VPWR _08974_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A VGND VGND VPWR VPWR _08831_/X sky130_fd_sc_hd__buf_1
XFILLER_112_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08762_/A _10133_/A VGND VGND VPWR VPWR _08762_/Y sky130_fd_sc_hd__nor2_1
X_08693_ _08876_/A _08691_/X _08876_/B VGND VGND VPWR VPWR _08693_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09314_ _09274_/A _09274_/B _09274_/X _10543_/A VGND VGND VPWR VPWR _10664_/A sky130_fd_sc_hd__a22o_1
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09245_ _08572_/A _09858_/A _09317_/A VGND VGND VPWR VPWR _09245_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09176_ _09175_/Y _09040_/Y _09143_/Y VGND VGND VPWR VPWR _09180_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10020_ _08844_/A _09070_/A _08944_/X _10019_/X VGND VGND VPWR VPWR _10020_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11971_ _11954_/Y _11969_/X _11970_/Y VGND VGND VPWR VPWR _11971_/X sky130_fd_sc_hd__o21a_1
XFILLER_17_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10922_ _14614_/A _10922_/B VGND VGND VPWR VPWR _10922_/X sky130_fd_sc_hd__or2_1
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13710_ _15046_/A _13503_/B _13503_/Y VGND VGND VPWR VPWR _13710_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14690_ _15347_/A _14661_/B _14661_/Y VGND VGND VPWR VPWR _14690_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10853_ _11942_/A _10708_/B _10708_/Y VGND VGND VPWR VPWR _10853_/Y sky130_fd_sc_hd__o21ai_1
X_13641_ _15122_/A _13641_/B VGND VGND VPWR VPWR _13641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16360_ _16329_/X _16359_/Y _16329_/X _16359_/Y VGND VGND VPWR VPWR _16407_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _12137_/A _12915_/B _12917_/A _12915_/Y VGND VGND VPWR VPWR _13572_/X sky130_fd_sc_hd__o2bb2a_1
X_10784_ _11980_/A _10784_/B VGND VGND VPWR VPWR _10784_/Y sky130_fd_sc_hd__nor2_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16291_ _16264_/A _16330_/A _16264_/Y VGND VGND VPWR VPWR _16291_/Y sky130_fd_sc_hd__o21ai_1
X_12523_ _13441_/A _11372_/B _11372_/Y VGND VGND VPWR VPWR _12524_/B sky130_fd_sc_hd__o21a_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15311_ _15341_/A _15341_/B VGND VGND VPWR VPWR _15375_/A sky130_fd_sc_hd__and2_1
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15242_ _15225_/X _15241_/Y _15225_/X _15241_/Y VGND VGND VPWR VPWR _15243_/B sky130_fd_sc_hd__a2bb2o_1
X_12454_ _12454_/A _12454_/B VGND VGND VPWR VPWR _12454_/Y sky130_fd_sc_hd__nor2_1
X_11405_ _11411_/B _11405_/B VGND VGND VPWR VPWR _12331_/A sky130_fd_sc_hd__or2_1
X_15173_ _15159_/Y _15172_/Y _15159_/Y _15172_/Y VGND VGND VPWR VPWR _15556_/B sky130_fd_sc_hd__a2bb2o_1
X_12385_ _12437_/A _12385_/B VGND VGND VPWR VPWR _12385_/Y sky130_fd_sc_hd__nor2_1
X_14124_ _14125_/A _14126_/A VGND VGND VPWR VPWR _14124_/Y sky130_fd_sc_hd__nor2_1
X_11336_ _11509_/A _11510_/B _11509_/A _11510_/B VGND VGND VPWR VPWR _11336_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14055_ _14055_/A _14055_/B VGND VGND VPWR VPWR _14055_/X sky130_fd_sc_hd__or2_1
XFILLER_106_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11267_ _13370_/A VGND VGND VPWR VPWR _14008_/A sky130_fd_sc_hd__inv_2
X_13006_ _15146_/A _12922_/B _12922_/Y VGND VGND VPWR VPWR _13006_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11198_ _09424_/A _09131_/B _09131_/Y VGND VGND VPWR VPWR _11199_/A sky130_fd_sc_hd__o21ai_1
X_10218_ _10216_/X _10217_/Y _10216_/X _10217_/Y VGND VGND VPWR VPWR _11232_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_121_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10149_ _10151_/A VGND VGND VPWR VPWR _10241_/B sky130_fd_sc_hd__buf_1
XFILLER_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14957_ _14956_/A _14956_/B _14956_/Y VGND VGND VPWR VPWR _14957_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14888_ _14820_/X _14887_/X _14820_/X _14887_/X VGND VGND VPWR VPWR _14914_/B sky130_fd_sc_hd__a2bb2o_1
X_13908_ _15410_/A _13951_/B VGND VGND VPWR VPWR _13908_/Y sky130_fd_sc_hd__nor2_1
X_13839_ _14645_/A _13839_/B VGND VGND VPWR VPWR _13839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15509_ _15509_/A _15509_/B VGND VGND VPWR VPWR _15510_/A sky130_fd_sc_hd__nand2_1
X_09030_ _09539_/B _09030_/B VGND VGND VPWR VPWR _09031_/B sky130_fd_sc_hd__or2_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09932_ _09932_/A _09932_/B VGND VGND VPWR VPWR _09932_/X sky130_fd_sc_hd__or2_1
XFILLER_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09863_ _09863_/A _09863_/B VGND VGND VPWR VPWR _09863_/X sky130_fd_sc_hd__or2_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08814_ _08814_/A VGND VGND VPWR VPWR _08814_/X sky130_fd_sc_hd__buf_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09794_/A VGND VGND VPWR VPWR _09794_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08745_ _08745_/A VGND VGND VPWR VPWR _08745_/Y sky130_fd_sc_hd__inv_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08676_ _10098_/B VGND VGND VPWR VPWR _08677_/B sky130_fd_sc_hd__inv_2
XFILLER_26_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09228_ _09228_/A _09228_/B VGND VGND VPWR VPWR _09800_/A sky130_fd_sc_hd__or2_1
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09159_ _08709_/Y _09158_/Y _08743_/X VGND VGND VPWR VPWR _09160_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12170_ _12170_/A VGND VGND VPWR VPWR _12170_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11121_ _12256_/A VGND VGND VPWR VPWR _13719_/A sky130_fd_sc_hd__buf_1
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11052_ _12039_/A _10894_/B _10894_/Y VGND VGND VPWR VPWR _11052_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15860_ _15860_/A VGND VGND VPWR VPWR _15900_/A sky130_fd_sc_hd__inv_2
XFILLER_88_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10003_ _10001_/X _10002_/X _10001_/X _10002_/X VGND VGND VPWR VPWR _10344_/B sky130_fd_sc_hd__o2bb2a_4
X_14811_ _14722_/X _14810_/X _14722_/X _14810_/X VGND VGND VPWR VPWR _14812_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15791_ _15787_/Y _15789_/Y _15790_/Y VGND VGND VPWR VPWR _15795_/B sky130_fd_sc_hd__o21ai_2
XFILLER_64_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14742_ _15349_/A _14742_/B VGND VGND VPWR VPWR _14742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11954_ _13083_/A _11970_/B VGND VGND VPWR VPWR _11954_/Y sky130_fd_sc_hd__nor2_1
X_10905_ _10767_/X _10904_/X _10767_/X _10904_/X VGND VGND VPWR VPWR _10910_/B sky130_fd_sc_hd__a2bb2o_1
X_11885_ _11885_/A _11898_/B VGND VGND VPWR VPWR _11885_/Y sky130_fd_sc_hd__nor2_1
X_14673_ _14673_/A _14673_/B VGND VGND VPWR VPWR _14673_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16412_ _16469_/Q VGND VGND VPWR VPWR _16412_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13624_ _13624_/A VGND VGND VPWR VPWR _15134_/A sky130_fd_sc_hd__buf_1
X_10836_ _10805_/X _10835_/X _10805_/X _10835_/X VGND VGND VPWR VPWR _10953_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16343_ _16343_/A VGND VGND VPWR VPWR _16343_/X sky130_fd_sc_hd__buf_1
X_10767_ _11063_/A _11065_/B VGND VGND VPWR VPWR _10767_/X sky130_fd_sc_hd__or2_1
X_13555_ _13555_/A _13555_/B VGND VGND VPWR VPWR _13556_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16274_ _16145_/Y _16271_/X _16273_/Y VGND VGND VPWR VPWR _16274_/Y sky130_fd_sc_hd__o21ai_1
X_12506_ _14137_/A VGND VGND VPWR VPWR _13445_/A sky130_fd_sc_hd__buf_1
X_10698_ _13512_/A _10804_/B _13512_/A _10804_/B VGND VGND VPWR VPWR _10698_/X sky130_fd_sc_hd__a2bb2o_1
X_13486_ _10673_/Y _11862_/A _10574_/Y _13485_/X VGND VGND VPWR VPWR _13486_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15225_ _15190_/A _15190_/B _15190_/Y _15224_/X VGND VGND VPWR VPWR _15225_/X sky130_fd_sc_hd__a2bb2o_1
X_12437_ _12437_/A _12437_/B VGND VGND VPWR VPWR _12437_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15156_ _15119_/A _15119_/B _15119_/Y _15155_/X VGND VGND VPWR VPWR _15156_/X sky130_fd_sc_hd__a2bb2o_1
X_14107_ _14107_/A _14111_/B VGND VGND VPWR VPWR _14107_/Y sky130_fd_sc_hd__nor2_1
X_12368_ _12367_/Y _12260_/X _12283_/Y VGND VGND VPWR VPWR _12368_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12299_ _14008_/A _12299_/B VGND VGND VPWR VPWR _12299_/Y sky130_fd_sc_hd__nand2_1
X_15087_ _15087_/A _15087_/B VGND VGND VPWR VPWR _15087_/X sky130_fd_sc_hd__or2_1
X_11319_ _10084_/X _11318_/X _10084_/X _11318_/X VGND VGND VPWR VPWR _11320_/B sky130_fd_sc_hd__a2bb2o_1
X_14038_ _14038_/A _14038_/B VGND VGND VPWR VPWR _14038_/X sky130_fd_sc_hd__and2_1
XFILLER_79_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15989_ _15973_/X _15988_/Y _15973_/X _15988_/Y VGND VGND VPWR VPWR _15991_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08530_ _09527_/A VGND VGND VPWR VPWR _09474_/B sky130_fd_sc_hd__inv_2
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08461_ _08460_/A _08308_/Y _08460_/Y _08308_/A _08441_/X VGND VGND VPWR VPWR _08697_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08392_ _08392_/A VGND VGND VPWR VPWR _08392_/Y sky130_fd_sc_hd__inv_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09013_ _08893_/X _09021_/S _08579_/Y VGND VGND VPWR VPWR _09020_/S sky130_fd_sc_hd__o21ai_1
XFILLER_105_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09915_ _09859_/A _09859_/B _09914_/Y VGND VGND VPWR VPWR _10948_/A sky130_fd_sc_hd__a21oi_1
XFILLER_98_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09846_ _10490_/B _10489_/A VGND VGND VPWR VPWR _09847_/B sky130_fd_sc_hd__or2_1
XFILLER_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09777_ _10079_/A _09775_/Y _09776_/Y VGND VGND VPWR VPWR _09779_/B sky130_fd_sc_hd__o21ai_1
XFILLER_85_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08728_ _08715_/A _08715_/B _08715_/X _08727_/X VGND VGND VPWR VPWR _08729_/A sky130_fd_sc_hd__a22o_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08659_ _10099_/B VGND VGND VPWR VPWR _08679_/B sky130_fd_sc_hd__buf_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _13132_/A VGND VGND VPWR VPWR _15433_/A sky130_fd_sc_hd__buf_1
XFILLER_53_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10621_ _10621_/A _12606_/A VGND VGND VPWR VPWR _15212_/A sky130_fd_sc_hd__or2_1
X_13340_ _13340_/A _13340_/B VGND VGND VPWR VPWR _13340_/X sky130_fd_sc_hd__and2_1
X_10552_ _10554_/A VGND VGND VPWR VPWR _10552_/Y sky130_fd_sc_hd__inv_2
X_13271_ _12045_/A _13270_/Y _12045_/A _13270_/Y VGND VGND VPWR VPWR _13272_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12222_ _12144_/X _12221_/X _12144_/X _12221_/X VGND VGND VPWR VPWR _12223_/B sky130_fd_sc_hd__a2bb2o_1
X_15010_ _15044_/A _15044_/B VGND VGND VPWR VPWR _15058_/A sky130_fd_sc_hd__and2_1
XFILLER_6_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10483_ _09849_/Y _10482_/X _09848_/X _09851_/B _10794_/A VGND VGND VPWR VPWR _12932_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12153_ _13901_/A _12153_/B VGND VGND VPWR VPWR _12153_/X sky130_fd_sc_hd__or2_1
XFILLER_78_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11104_ _11006_/A _10926_/X _11005_/X VGND VGND VPWR VPWR _11104_/X sky130_fd_sc_hd__o21a_1
X_12084_ _12084_/A _12084_/B VGND VGND VPWR VPWR _12084_/Y sky130_fd_sc_hd__nor2_1
X_15912_ _15978_/A _15978_/B VGND VGND VPWR VPWR _15912_/Y sky130_fd_sc_hd__nand2_1
X_11035_ _13913_/A _11086_/B VGND VGND VPWR VPWR _11217_/A sky130_fd_sc_hd__and2_1
XFILLER_89_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15843_ _14219_/A _15842_/X _12622_/X VGND VGND VPWR VPWR _15843_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15774_ _12611_/A _15773_/A _12611_/Y _15773_/Y VGND VGND VPWR VPWR _15775_/B sky130_fd_sc_hd__o22a_1
X_12986_ _12933_/X _12985_/Y _12933_/X _12985_/Y VGND VGND VPWR VPWR _13021_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14725_ _14807_/A _14723_/X _14807_/B VGND VGND VPWR VPWR _14725_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11937_ _11936_/A _11983_/B _11936_/Y VGND VGND VPWR VPWR _11937_/Y sky130_fd_sc_hd__o21ai_1
X_14656_ _14621_/Y _14654_/X _14655_/Y VGND VGND VPWR VPWR _14656_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11868_ _10545_/X _11914_/B _10545_/X _11914_/B VGND VGND VPWR VPWR _11868_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14587_ _14587_/A _14587_/B VGND VGND VPWR VPWR _14587_/Y sky130_fd_sc_hd__nand2_1
X_13607_ _13572_/X _13606_/Y _13572_/X _13606_/Y VGND VGND VPWR VPWR _13608_/B sky130_fd_sc_hd__a2bb2o_1
X_11799_ _13563_/A _11778_/B _11778_/X _11798_/X VGND VGND VPWR VPWR _11799_/X sky130_fd_sc_hd__o22a_1
X_10819_ _10819_/A VGND VGND VPWR VPWR _12084_/A sky130_fd_sc_hd__inv_2
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16326_ _16326_/A _16326_/B VGND VGND VPWR VPWR _16326_/Y sky130_fd_sc_hd__nand2_1
X_13538_ _15042_/A _13509_/B _13509_/Y _13537_/X VGND VGND VPWR VPWR _13538_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16257_ _16257_/A VGND VGND VPWR VPWR _16324_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13469_ _13465_/X _13468_/X _13465_/X _13468_/X VGND VGND VPWR VPWR _13469_/X sky130_fd_sc_hd__a2bb2o_1
X_16188_ _16105_/X _16187_/X _16105_/X _16187_/X VGND VGND VPWR VPWR _16189_/B sky130_fd_sc_hd__a2bb2oi_1
X_15208_ _15208_/A _15208_/B VGND VGND VPWR VPWR _15208_/Y sky130_fd_sc_hd__nand2_1
X_15139_ _15089_/X _15138_/Y _15089_/X _15138_/Y VGND VGND VPWR VPWR _15140_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09700_ _09700_/A VGND VGND VPWR VPWR _09700_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09631_ _09952_/A _09631_/B VGND VGND VPWR VPWR _09632_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09562_ _09567_/A _09560_/X _09567_/B VGND VGND VPWR VPWR _09562_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08513_ _09863_/A _08509_/A _08464_/A _08512_/X _08464_/Y VGND VGND VPWR VPWR _08989_/A
+ sky130_fd_sc_hd__a32o_1
X_09493_ _08806_/A _09466_/X _08806_/A _09466_/X VGND VGND VPWR VPWR _09494_/B sky130_fd_sc_hd__o2bb2a_1
X_08444_ _08711_/A VGND VGND VPWR VPWR _09332_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08375_ input4/X _08248_/B _08317_/B _08447_/A VGND VGND VPWR VPWR _08375_/X sky130_fd_sc_hd__o22a_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09829_ _09829_/A _09829_/B VGND VGND VPWR VPWR _09830_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12840_ _12826_/Y _12838_/X _12839_/Y VGND VGND VPWR VPWR _12840_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12771_ _12751_/Y _12769_/X _12770_/Y VGND VGND VPWR VPWR _12771_/X sky130_fd_sc_hd__o21a_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15485_/X _15489_/X _15485_/X _15489_/X VGND VGND VPWR VPWR _15552_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _14564_/A _14508_/X _14509_/X VGND VGND VPWR VPWR _14510_/X sky130_fd_sc_hd__o21a_1
X_11722_ _11722_/A _11722_/B VGND VGND VPWR VPWR _11722_/Y sky130_fd_sc_hd__nor2_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11652_/Y _11488_/Y _11552_/Y VGND VGND VPWR VPWR _11653_/X sky130_fd_sc_hd__o21a_1
X_14441_ _14468_/A _14468_/B VGND VGND VPWR VPWR _14441_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14372_ _14372_/A VGND VGND VPWR VPWR _14372_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10604_ _10604_/A VGND VGND VPWR VPWR _10604_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16111_ _16073_/X _16109_/X _16171_/B VGND VGND VPWR VPWR _16111_/X sky130_fd_sc_hd__o21a_1
X_13323_ _14736_/A _13294_/B _13294_/Y VGND VGND VPWR VPWR _13323_/Y sky130_fd_sc_hd__o21ai_1
X_11584_ _09169_/A _09362_/A _09429_/X VGND VGND VPWR VPWR _11584_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10535_ _09898_/A _09898_/B _09898_/X VGND VGND VPWR VPWR _10535_/X sky130_fd_sc_hd__o21ba_1
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16042_ _16042_/A _16042_/B VGND VGND VPWR VPWR _16042_/Y sky130_fd_sc_hd__nand2_1
X_13254_ _13189_/X _13253_/Y _13189_/X _13253_/Y VGND VGND VPWR VPWR _13282_/B sky130_fd_sc_hd__a2bb2o_1
X_10466_ _10466_/A VGND VGND VPWR VPWR _10466_/Y sky130_fd_sc_hd__clkinvlp_2
X_12205_ _14011_/A _12205_/B VGND VGND VPWR VPWR _12205_/Y sky130_fd_sc_hd__nand2_1
X_13185_ _13178_/Y _13183_/X _13184_/Y VGND VGND VPWR VPWR _13185_/X sky130_fd_sc_hd__o21a_1
X_12136_ _12137_/A _12137_/B VGND VGND VPWR VPWR _12136_/X sky130_fd_sc_hd__or2_1
X_10397_ _11778_/A VGND VGND VPWR VPWR _13563_/A sky130_fd_sc_hd__buf_1
XFILLER_96_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12067_ _12106_/A VGND VGND VPWR VPWR _13200_/A sky130_fd_sc_hd__buf_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11018_ _12851_/A VGND VGND VPWR VPWR _15066_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15826_ _15697_/X _15825_/Y _15703_/Y VGND VGND VPWR VPWR _15826_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15757_ _14911_/X _15756_/X _14911_/X _15756_/X VGND VGND VPWR VPWR _15758_/B sky130_fd_sc_hd__a2bb2oi_1
X_12969_ _14599_/A _12942_/B _12942_/Y VGND VGND VPWR VPWR _12969_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15688_ _14399_/Y _15687_/Y _14399_/Y _15687_/Y VGND VGND VPWR VPWR _15694_/B sky130_fd_sc_hd__a2bb2o_1
X_14708_ _15335_/A _14649_/B _14649_/Y VGND VGND VPWR VPWR _14708_/Y sky130_fd_sc_hd__o21ai_1
X_14639_ _14572_/X _14638_/Y _14572_/X _14638_/Y VGND VGND VPWR VPWR _14645_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16309_ _16251_/A _16318_/A _16251_/Y VGND VGND VPWR VPWR _16309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08993_ _09340_/A _08748_/Y _09341_/A VGND VGND VPWR VPWR _08993_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09614_ _09548_/X _09613_/Y _09548_/X _09613_/Y VGND VGND VPWR VPWR _09652_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09545_ _09538_/A _09538_/B _09538_/X _09544_/X VGND VGND VPWR VPWR _09546_/A sky130_fd_sc_hd__o22a_1
XFILLER_36_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09476_ _10009_/A _09476_/B VGND VGND VPWR VPWR _09476_/X sky130_fd_sc_hd__or2_1
XFILLER_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08427_ _08714_/A VGND VGND VPWR VPWR _08794_/A sky130_fd_sc_hd__buf_1
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08358_ _08358_/A input18/X VGND VGND VPWR VPWR _08399_/A sky130_fd_sc_hd__nor2_1
X_08289_ _08336_/A input31/X _08337_/A _08339_/A VGND VGND VPWR VPWR _08334_/A sky130_fd_sc_hd__o22a_1
XFILLER_118_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10320_ _09958_/A _09958_/B _09958_/Y VGND VGND VPWR VPWR _10320_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10251_ _10251_/A VGND VGND VPWR VPWR _10251_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10182_ _10182_/A VGND VGND VPWR VPWR _10182_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14990_ _12433_/X _14989_/X _12433_/X _14989_/X VGND VGND VPWR VPWR _14990_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_115_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13941_ _15400_/A _13941_/B VGND VGND VPWR VPWR _13941_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13872_ _13872_/A _13872_/B VGND VGND VPWR VPWR _13873_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15611_ _16040_/A VGND VGND VPWR VPWR _15677_/A sky130_fd_sc_hd__inv_2
XFILLER_74_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12823_ _12841_/A _12841_/B VGND VGND VPWR VPWR _12823_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15542_ _15542_/A _15542_/B VGND VGND VPWR VPWR _15542_/X sky130_fd_sc_hd__or2_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12768_/A _12768_/B VGND VGND VPWR VPWR _12754_/Y sky130_fd_sc_hd__nor2_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11699_/X _11704_/Y _11699_/X _11704_/Y VGND VGND VPWR VPWR _11705_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15473_ _15473_/A _15473_/B VGND VGND VPWR VPWR _15473_/Y sky130_fd_sc_hd__nand2_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12685_/A _12685_/B VGND VGND VPWR VPWR _12685_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14424_ _14424_/A _14424_/B VGND VGND VPWR VPWR _14424_/Y sky130_fd_sc_hd__nor2_1
X_11636_ _11634_/Y _11635_/Y _11543_/Y VGND VGND VPWR VPWR _11636_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14355_ _14249_/Y _14354_/Y _14249_/Y _14354_/Y VGND VGND VPWR VPWR _14377_/A sky130_fd_sc_hd__a2bb2o_1
X_11567_ _12410_/A _11567_/B VGND VGND VPWR VPWR _11567_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14286_ _14282_/X _14284_/X _14398_/B VGND VGND VPWR VPWR _14286_/X sky130_fd_sc_hd__o21a_1
X_13306_ _14858_/A _13306_/B VGND VGND VPWR VPWR _13306_/Y sky130_fd_sc_hd__nand2_1
X_10518_ _11794_/A _10429_/B _11794_/A _10429_/B VGND VGND VPWR VPWR _10518_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16025_ _16030_/A _16030_/B VGND VGND VPWR VPWR _16025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13237_ _14473_/A VGND VGND VPWR VPWR _14734_/A sky130_fd_sc_hd__buf_1
XFILLER_7_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11498_ _11593_/A _11498_/B VGND VGND VPWR VPWR _12393_/A sky130_fd_sc_hd__or2_2
X_10449_ _11806_/A VGND VGND VPWR VPWR _11767_/A sky130_fd_sc_hd__inv_2
XFILLER_130_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13168_ _13190_/A _13190_/B VGND VGND VPWR VPWR _13168_/Y sky130_fd_sc_hd__nor2_1
X_13099_ _13009_/A _13098_/Y _13009_/A _13098_/Y VGND VGND VPWR VPWR _13101_/B sky130_fd_sc_hd__a2bb2o_1
X_12119_ _13192_/A _12059_/B _12059_/Y VGND VGND VPWR VPWR _12119_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15809_ _16108_/A _15809_/B VGND VGND VPWR VPWR _15809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09330_ _09330_/A _09330_/B VGND VGND VPWR VPWR _10035_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09261_ _10242_/A VGND VGND VPWR VPWR _09262_/B sky130_fd_sc_hd__buf_1
XFILLER_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09192_ _09561_/B _09156_/X _09190_/Y _11667_/B VGND VGND VPWR VPWR _09193_/A sky130_fd_sc_hd__o22a_1
XFILLER_119_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08976_ _08976_/A _08976_/B VGND VGND VPWR VPWR _11373_/B sky130_fd_sc_hd__or2_1
XFILLER_84_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09528_ _09528_/A VGND VGND VPWR VPWR _09528_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09459_ _09459_/A _09459_/B VGND VGND VPWR VPWR _09459_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12470_ _12439_/X _12469_/X _12439_/X _12469_/X VGND VGND VPWR VPWR _12470_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11421_ _13404_/A _11422_/B VGND VGND VPWR VPWR _12607_/B sky130_fd_sc_hd__or2_1
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14140_ _14140_/A _14065_/X VGND VGND VPWR VPWR _14140_/X sky130_fd_sc_hd__or2b_1
X_11352_ _13889_/A _11352_/B VGND VGND VPWR VPWR _11352_/X sky130_fd_sc_hd__or2_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10303_ _10303_/A VGND VGND VPWR VPWR _11762_/A sky130_fd_sc_hd__inv_4
X_14071_ _14069_/X _14070_/X _14069_/X _14070_/X VGND VGND VPWR VPWR _14071_/X sky130_fd_sc_hd__a2bb2o_1
X_11283_ _11586_/A _11283_/B VGND VGND VPWR VPWR _12292_/A sky130_fd_sc_hd__or2_2
XFILLER_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13022_ _13075_/A _13020_/X _13021_/X VGND VGND VPWR VPWR _13022_/X sky130_fd_sc_hd__o21a_1
X_10234_ _10234_/A VGND VGND VPWR VPWR _10234_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10165_ _10167_/A VGND VGND VPWR VPWR _10468_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14973_ _12431_/A _12424_/Y _14973_/B1 _14936_/X VGND VGND VPWR VPWR _14973_/Y sky130_fd_sc_hd__o22ai_2
X_10096_ _10215_/A _11239_/A VGND VGND VPWR VPWR _11736_/A sky130_fd_sc_hd__or2_1
X_13924_ _15402_/A _13943_/B VGND VGND VPWR VPWR _13924_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13855_ _14409_/A _13855_/B VGND VGND VPWR VPWR _13855_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12806_ _12776_/A _12776_/B _12776_/Y VGND VGND VPWR VPWR _12806_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10998_ _13702_/A _11115_/B _10997_/Y VGND VGND VPWR VPWR _10998_/Y sky130_fd_sc_hd__o21ai_1
X_13786_ _12859_/A _13785_/B _13867_/A VGND VGND VPWR VPWR _13786_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15525_ _15521_/Y _15632_/A _15524_/Y VGND VGND VPWR VPWR _15529_/B sky130_fd_sc_hd__o21ai_1
XFILLER_70_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12691_/A _12691_/B _12691_/Y VGND VGND VPWR VPWR _12737_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15456_ _15456_/A _15406_/X VGND VGND VPWR VPWR _15456_/X sky130_fd_sc_hd__or2b_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _10814_/Y _12667_/Y _10687_/Y VGND VGND VPWR VPWR _12669_/A sky130_fd_sc_hd__o21ai_1
X_14407_ _14407_/A VGND VGND VPWR VPWR _15552_/A sky130_fd_sc_hd__buf_1
X_11619_ _11619_/A _11619_/B VGND VGND VPWR VPWR _11619_/Y sky130_fd_sc_hd__nor2_1
X_12599_ _12599_/A VGND VGND VPWR VPWR _12599_/Y sky130_fd_sc_hd__clkinvlp_2
X_15387_ _15387_/A _15333_/X VGND VGND VPWR VPWR _15387_/X sky130_fd_sc_hd__or2b_1
XFILLER_128_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14338_ _14100_/A _13425_/B _13425_/Y VGND VGND VPWR VPWR _14338_/X sky130_fd_sc_hd__o21a_1
X_14269_ _14197_/Y _14267_/Y _14268_/Y VGND VGND VPWR VPWR _14270_/A sky130_fd_sc_hd__o21ai_2
X_16008_ _15930_/X _16008_/B VGND VGND VPWR VPWR _16008_/Y sky130_fd_sc_hd__nand2b_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08830_/A VGND VGND VPWR VPWR _08831_/A sky130_fd_sc_hd__inv_2
XFILLER_112_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _10009_/A VGND VGND VPWR VPWR _08762_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08692_ _08692_/A _10119_/B VGND VGND VPWR VPWR _08876_/B sky130_fd_sc_hd__and2_1
XFILLER_53_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09313_ _10437_/A _09311_/Y _09312_/Y VGND VGND VPWR VPWR _10543_/A sky130_fd_sc_hd__o21ai_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09244_ _09555_/A _09734_/A VGND VGND VPWR VPWR _09317_/A sky130_fd_sc_hd__or2_1
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09175_ _09432_/A _09175_/B VGND VGND VPWR VPWR _09175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08959_ _08681_/Y _08958_/X _08681_/Y _08958_/X VGND VGND VPWR VPWR _11399_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11970_ _11970_/A _11970_/B VGND VGND VPWR VPWR _11970_/Y sky130_fd_sc_hd__nand2_1
X_10921_ _10921_/A VGND VGND VPWR VPWR _14614_/A sky130_fd_sc_hd__buf_1
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10852_ _12063_/A VGND VGND VPWR VPWR _10921_/A sky130_fd_sc_hd__inv_2
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13640_ _13640_/A VGND VGND VPWR VPWR _15122_/A sky130_fd_sc_hd__buf_1
XFILLER_32_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10783_ _13058_/A VGND VGND VPWR VPWR _12068_/A sky130_fd_sc_hd__buf_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _14428_/A _13573_/B VGND VGND VPWR VPWR _13571_/X sky130_fd_sc_hd__and2_1
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16290_ _16332_/A _16332_/B VGND VGND VPWR VPWR _16290_/Y sky130_fd_sc_hd__nor2_1
X_12522_ _14125_/A VGND VGND VPWR VPWR _13441_/A sky130_fd_sc_hd__buf_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15310_ _15277_/X _15309_/Y _15277_/X _15309_/Y VGND VGND VPWR VPWR _15341_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15241_ _15187_/A _15187_/B _15187_/Y VGND VGND VPWR VPWR _15241_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12453_ _12450_/X _12452_/X _12450_/X _12452_/X VGND VGND VPWR VPWR _12454_/B sky130_fd_sc_hd__a2bb2o_1
X_15172_ _15171_/A _15425_/B _15171_/Y VGND VGND VPWR VPWR _15172_/Y sky130_fd_sc_hd__o21ai_1
X_12384_ _12420_/B _12383_/Y _12420_/B _12383_/Y VGND VGND VPWR VPWR _12385_/B sky130_fd_sc_hd__a2bb2o_1
X_11404_ _08951_/Y _11403_/X _08951_/Y _11403_/X VGND VGND VPWR VPWR _11405_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14123_ _14058_/X _14122_/X _14058_/X _14122_/X VGND VGND VPWR VPWR _14126_/A sky130_fd_sc_hd__a2bb2o_1
X_11335_ _11315_/X _11334_/X _11315_/X _11334_/X VGND VGND VPWR VPWR _11510_/B sky130_fd_sc_hd__a2bb2o_1
X_14054_ _14108_/A _14023_/B _14023_/X _14053_/X VGND VGND VPWR VPWR _14054_/X sky130_fd_sc_hd__o22a_1
X_11266_ _09179_/Y _11265_/A _09179_/A _11265_/Y _09204_/X VGND VGND VPWR VPWR _13370_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13005_ _13005_/A VGND VGND VPWR VPWR _15146_/A sky130_fd_sc_hd__buf_1
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10217_ _10059_/A _10059_/B _10059_/Y VGND VGND VPWR VPWR _10217_/Y sky130_fd_sc_hd__a21oi_1
X_11197_ _14057_/A _11197_/B VGND VGND VPWR VPWR _11197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10148_ _10117_/A _10117_/B _10118_/A VGND VGND VPWR VPWR _10151_/A sky130_fd_sc_hd__a21bo_1
X_14956_ _14956_/A _14956_/B VGND VGND VPWR VPWR _14956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10079_ _10079_/A _10079_/B VGND VGND VPWR VPWR _10816_/B sky130_fd_sc_hd__or2_1
X_13907_ _13850_/X _13906_/Y _13850_/X _13906_/Y VGND VGND VPWR VPWR _13951_/B sky130_fd_sc_hd__a2bb2o_1
X_14887_ _14798_/A _14798_/B _14798_/A _14798_/B VGND VGND VPWR VPWR _14887_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13838_ _10909_/A _13836_/Y _13837_/Y VGND VGND VPWR VPWR _13838_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13769_ _13809_/A _13767_/X _13768_/X VGND VGND VPWR VPWR _13769_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15508_ _12237_/X _15507_/Y _12237_/X _15507_/Y VGND VGND VPWR VPWR _15509_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15439_ _15417_/X _15438_/Y _15417_/X _15438_/Y VGND VGND VPWR VPWR _15440_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09931_ _09928_/X _09931_/B VGND VGND VPWR VPWR _09932_/B sky130_fd_sc_hd__nand2b_1
XFILLER_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09862_ _09862_/A _09924_/A VGND VGND VPWR VPWR _09863_/B sky130_fd_sc_hd__or2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08813_ _08813_/A VGND VGND VPWR VPWR _08814_/A sky130_fd_sc_hd__inv_2
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09793_/A _09793_/B VGND VGND VPWR VPWR _09794_/A sky130_fd_sc_hd__or2_1
XFILLER_100_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08744_ _08709_/Y _08742_/Y _08743_/X VGND VGND VPWR VPWR _08745_/A sky130_fd_sc_hd__o21ai_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08675_ _08664_/X _08402_/X _10228_/A _08674_/Y VGND VGND VPWR VPWR _10098_/B sky130_fd_sc_hd__a31o_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09227_ _09458_/B _09690_/A VGND VGND VPWR VPWR _09227_/X sky130_fd_sc_hd__or2_1
XFILLER_108_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09158_ _09158_/A VGND VGND VPWR VPWR _09158_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09089_ _10015_/B _09074_/B _09075_/B VGND VGND VPWR VPWR _09701_/A sky130_fd_sc_hd__a21bo_1
XFILLER_107_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11120_ _09966_/Y _11119_/A _10083_/A _11119_/Y _11593_/A VGND VGND VPWR VPWR _12256_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11051_ _12141_/A VGND VGND VPWR VPWR _13925_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10002_ _09521_/Y _09792_/A _09521_/Y _09792_/A VGND VGND VPWR VPWR _10002_/X sky130_fd_sc_hd__o2bb2a_1
X_14810_ _15398_/A _14717_/B _15398_/A _14717_/B VGND VGND VPWR VPWR _14810_/X sky130_fd_sc_hd__a2bb2o_1
X_15790_ _16089_/A _15790_/B VGND VGND VPWR VPWR _15790_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14741_ _14776_/A _14739_/X _14740_/X VGND VGND VPWR VPWR _14741_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11953_ _11900_/A _11952_/Y _11900_/A _11952_/Y VGND VGND VPWR VPWR _11970_/B sky130_fd_sc_hd__a2bb2o_1
X_10904_ _10904_/A _10769_/X VGND VGND VPWR VPWR _10904_/X sky130_fd_sc_hd__or2b_1
X_11884_ _11839_/X _11883_/Y _11839_/X _11883_/Y VGND VGND VPWR VPWR _11898_/B sky130_fd_sc_hd__a2bb2o_1
X_14672_ _12185_/Y _14671_/X _12185_/Y _14671_/X VGND VGND VPWR VPWR _14673_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16411_ _16454_/A _16411_/B VGND VGND VPWR VPWR _16474_/D sky130_fd_sc_hd__or2_1
X_13623_ _13623_/A VGND VGND VPWR VPWR _13623_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10835_ _13509_/A _10955_/B _13509_/A _10955_/B VGND VGND VPWR VPWR _10835_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16342_ _16361_/A VGND VGND VPWR VPWR _16343_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10766_ _10766_/A _13008_/A VGND VGND VPWR VPWR _11065_/B sky130_fd_sc_hd__nand2_1
X_13554_ _13534_/X _13553_/Y _13534_/X _13553_/Y VGND VGND VPWR VPWR _13555_/B sky130_fd_sc_hd__a2bb2o_1
X_16273_ _16273_/A _16338_/A VGND VGND VPWR VPWR _16273_/Y sky130_fd_sc_hd__nand2_1
X_12505_ _12640_/A _12640_/B VGND VGND VPWR VPWR _14170_/A sky130_fd_sc_hd__and2_1
X_13485_ _10552_/Y _11813_/A _10474_/Y _13484_/X VGND VGND VPWR VPWR _13485_/X sky130_fd_sc_hd__o22a_1
X_10697_ _10676_/X _10696_/X _10676_/X _10696_/X VGND VGND VPWR VPWR _10804_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15224_ _15193_/A _15193_/B _15193_/Y _15223_/X VGND VGND VPWR VPWR _15224_/X sky130_fd_sc_hd__a2bb2o_1
X_12436_ _13494_/A _12435_/B _12435_/Y VGND VGND VPWR VPWR _12439_/A sky130_fd_sc_hd__a21oi_1
X_15155_ _15122_/A _15122_/B _15122_/Y _15154_/X VGND VGND VPWR VPWR _15155_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14106_ _14102_/Y _14104_/Y _14105_/Y VGND VGND VPWR VPWR _14111_/B sky130_fd_sc_hd__o21ai_2
XFILLER_99_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12367_ _13788_/A _12367_/B VGND VGND VPWR VPWR _12367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12298_ _12250_/X _12297_/Y _12250_/X _12297_/Y VGND VGND VPWR VPWR _12299_/B sky130_fd_sc_hd__a2bb2o_1
X_15086_ _15087_/A _15087_/B VGND VGND VPWR VPWR _15144_/A sky130_fd_sc_hd__and2_1
X_11318_ _10040_/X _11318_/B VGND VGND VPWR VPWR _11318_/X sky130_fd_sc_hd__and2b_1
X_11249_ _11247_/X _11248_/X _11247_/X _11248_/X VGND VGND VPWR VPWR _11252_/B sky130_fd_sc_hd__a2bb2o_1
X_14037_ _13940_/Y _14036_/X _13940_/Y _14036_/X VGND VGND VPWR VPWR _14038_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15988_ _15981_/X _15988_/B VGND VGND VPWR VPWR _15988_/Y sky130_fd_sc_hd__nand2b_1
X_14939_ _14934_/A _14938_/B _14938_/Y VGND VGND VPWR VPWR _14939_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08460_ _08460_/A VGND VGND VPWR VPWR _08460_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08391_ input9/X _08279_/B _08279_/Y VGND VGND VPWR VPWR _08392_/A sky130_fd_sc_hd__a21oi_2
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09012_ _08795_/X _09011_/Y _09213_/B VGND VGND VPWR VPWR _09021_/S sky130_fd_sc_hd__a21oi_1
XFILLER_132_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09914_ _09914_/A VGND VGND VPWR VPWR _09914_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09845_ _09801_/A _09801_/B _09844_/Y VGND VGND VPWR VPWR _10489_/A sky130_fd_sc_hd__a21oi_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09776_ _09776_/A _09776_/B VGND VGND VPWR VPWR _09776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08727_ _08716_/A _08716_/B _08716_/X _08726_/X VGND VGND VPWR VPWR _08727_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08658_ _08657_/Y _08403_/Y _08657_/Y _08403_/Y VGND VGND VPWR VPWR _10099_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08589_ _08589_/A _08589_/B VGND VGND VPWR VPWR _09455_/B sky130_fd_sc_hd__or2_1
XFILLER_14_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10620_ _10522_/A _10619_/Y _10522_/A _10619_/Y VGND VGND VPWR VPWR _10629_/B sky130_fd_sc_hd__a2bb2o_1
X_10551_ _11853_/A VGND VGND VPWR VPWR _13515_/A sky130_fd_sc_hd__buf_1
XFILLER_127_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13270_ _15329_/A _13182_/B _13182_/Y VGND VGND VPWR VPWR _13270_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10482_ _09848_/A _09848_/B _09848_/X VGND VGND VPWR VPWR _10482_/X sky130_fd_sc_hd__o21ba_1
XFILLER_10_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12221_ _12221_/A _12145_/X VGND VGND VPWR VPWR _12221_/X sky130_fd_sc_hd__or2b_1
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12152_ _12212_/A _12150_/X _12151_/X VGND VGND VPWR VPWR _12152_/X sky130_fd_sc_hd__o21a_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11103_ _15057_/A VGND VGND VPWR VPWR _13893_/A sky130_fd_sc_hd__buf_1
X_12083_ _12082_/A _12082_/B _12082_/X _11999_/B VGND VGND VPWR VPWR _12174_/B sky130_fd_sc_hd__a22o_1
XFILLER_1_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15911_ _14170_/X _15851_/X _14170_/X _15851_/X VGND VGND VPWR VPWR _15978_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_104_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11034_ _10916_/X _11033_/X _10916_/X _11033_/X VGND VGND VPWR VPWR _11086_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15842_ _12594_/X _15841_/X _14225_/B VGND VGND VPWR VPWR _15842_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15773_ _15773_/A VGND VGND VPWR VPWR _15773_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12985_ _14466_/A _12934_/B _12934_/Y VGND VGND VPWR VPWR _12985_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14724_ _14724_/A _14724_/B VGND VGND VPWR VPWR _14807_/B sky130_fd_sc_hd__and2_1
X_11936_ _11936_/A _11983_/B VGND VGND VPWR VPWR _11936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14655_ _15341_/A _14655_/B VGND VGND VPWR VPWR _14655_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11867_ _11916_/B _11866_/Y _11916_/B _11866_/Y VGND VGND VPWR VPWR _11914_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14586_ _14542_/Y _14584_/X _14585_/Y VGND VGND VPWR VPWR _14586_/X sky130_fd_sc_hd__o21a_1
X_13606_ _13571_/X _13606_/B VGND VGND VPWR VPWR _13606_/Y sky130_fd_sc_hd__nand2b_1
X_11798_ _13567_/A _11783_/B _11783_/X _11797_/X VGND VGND VPWR VPWR _11798_/X sky130_fd_sc_hd__o22a_1
X_10818_ _10968_/A _10818_/B VGND VGND VPWR VPWR _10819_/A sky130_fd_sc_hd__or2_1
XFILLER_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16325_ _16302_/Y _16323_/X _16324_/Y VGND VGND VPWR VPWR _16325_/X sky130_fd_sc_hd__o21a_1
X_10749_ _13088_/A _10749_/B VGND VGND VPWR VPWR _10749_/Y sky130_fd_sc_hd__nand2_1
X_13537_ _15040_/A _13512_/B _13512_/Y _13536_/X VGND VGND VPWR VPWR _13537_/X sky130_fd_sc_hd__a2bb2o_1
X_16256_ _16211_/Y _16254_/X _16255_/Y VGND VGND VPWR VPWR _16256_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15207_ _15148_/X _15206_/Y _15148_/X _15206_/Y VGND VGND VPWR VPWR _15208_/B sky130_fd_sc_hd__a2bb2o_1
X_13468_ _13466_/Y _13467_/X _13466_/Y _13467_/X VGND VGND VPWR VPWR _13468_/X sky130_fd_sc_hd__a2bb2o_1
X_16187_ _16079_/X _16187_/B VGND VGND VPWR VPWR _16187_/X sky130_fd_sc_hd__and2b_1
X_13399_ _15519_/A VGND VGND VPWR VPWR _14090_/A sky130_fd_sc_hd__inv_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12419_ _12419_/A VGND VGND VPWR VPWR _12683_/A sky130_fd_sc_hd__buf_1
XFILLER_126_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15138_ _15081_/A _15081_/B _15081_/Y VGND VGND VPWR VPWR _15138_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15069_ _15069_/A _15069_/B VGND VGND VPWR VPWR _15069_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09630_ _09707_/A _09628_/Y _08929_/B _09629_/X VGND VGND VPWR VPWR _09631_/B sky130_fd_sc_hd__o22a_1
X_09561_ _09561_/A _09561_/B VGND VGND VPWR VPWR _09567_/B sky130_fd_sc_hd__and2_1
XFILLER_82_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08512_ _09345_/B _09791_/C VGND VGND VPWR VPWR _08512_/X sky130_fd_sc_hd__or2_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09492_ _09492_/A _09492_/B VGND VGND VPWR VPWR _09492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08443_ _08554_/A VGND VGND VPWR VPWR _08711_/A sky130_fd_sc_hd__inv_2
XFILLER_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08374_ input3/X _08251_/B _08322_/B _08440_/A VGND VGND VPWR VPWR _08447_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09828_ _10102_/A _09829_/A _09503_/B _09827_/X VGND VGND VPWR VPWR _09832_/A sky130_fd_sc_hd__a31o_1
XFILLER_104_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09759_ _10043_/A VGND VGND VPWR VPWR _10083_/A sky130_fd_sc_hd__buf_6
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12770_ _12770_/A _12770_/B VGND VGND VPWR VPWR _12770_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _12832_/A _11719_/A _10425_/A _11720_/Y VGND VGND VPWR VPWR _11722_/B sky130_fd_sc_hd__o22a_1
XFILLER_42_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11652_ _12396_/A _11652_/B VGND VGND VPWR VPWR _11652_/Y sky130_fd_sc_hd__nor2_1
X_14440_ _14435_/X _14439_/X _14435_/X _14439_/X VGND VGND VPWR VPWR _14468_/B sky130_fd_sc_hd__a2bb2o_1
X_14371_ _14371_/A _14371_/B VGND VGND VPWR VPWR _14372_/A sky130_fd_sc_hd__or2_1
XFILLER_23_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10603_ _09714_/A _09714_/B _09714_/Y VGND VGND VPWR VPWR _10604_/A sky130_fd_sc_hd__a21oi_1
XFILLER_127_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16110_ _16110_/A _16110_/B VGND VGND VPWR VPWR _16171_/B sky130_fd_sc_hd__or2_1
X_13322_ _13366_/A _13366_/B VGND VGND VPWR VPWR _13384_/A sky130_fd_sc_hd__and2_1
X_11583_ _11558_/A _11483_/X _11557_/X VGND VGND VPWR VPWR _11583_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10534_ _10481_/Y _10532_/X _10533_/Y VGND VGND VPWR VPWR _10534_/X sky130_fd_sc_hd__o21a_1
X_16041_ _16010_/Y _16039_/X _16040_/Y VGND VGND VPWR VPWR _16041_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13253_ _13190_/A _13190_/B _13190_/Y VGND VGND VPWR VPWR _13253_/Y sky130_fd_sc_hd__o21ai_1
X_10465_ _11857_/A _10556_/B _10464_/Y VGND VGND VPWR VPWR _10466_/A sky130_fd_sc_hd__o21ai_2
XFILLER_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12204_ _12156_/X _12203_/Y _12156_/X _12203_/Y VGND VGND VPWR VPWR _12205_/B sky130_fd_sc_hd__a2bb2o_1
X_13184_ _13184_/A _13184_/B VGND VGND VPWR VPWR _13184_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10396_ _10396_/A VGND VGND VPWR VPWR _11778_/A sky130_fd_sc_hd__buf_1
XFILLER_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12135_ _12044_/A _12134_/X _12044_/A _12134_/X VGND VGND VPWR VPWR _12137_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12066_ _12016_/Y _12064_/X _12065_/Y VGND VGND VPWR VPWR _12066_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11017_ _13547_/A VGND VGND VPWR VPWR _12851_/A sky130_fd_sc_hd__buf_1
X_15825_ _15991_/A _15825_/B VGND VGND VPWR VPWR _15825_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15756_ _14912_/A _14912_/B _14912_/Y VGND VGND VPWR VPWR _15756_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12968_ _13702_/A VGND VGND VPWR VPWR _14591_/A sky130_fd_sc_hd__inv_2
XFILLER_52_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15687_ _14397_/X _15687_/B VGND VGND VPWR VPWR _15687_/Y sky130_fd_sc_hd__nand2b_1
X_14707_ _14728_/A _14728_/B VGND VGND VPWR VPWR _14800_/A sky130_fd_sc_hd__and2_1
X_12899_ _12844_/X _12898_/Y _12844_/X _12898_/Y VGND VGND VPWR VPWR _12932_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11919_ _11919_/A VGND VGND VPWR VPWR _11987_/A sky130_fd_sc_hd__inv_2
X_14638_ _15272_/A _14573_/B _14573_/Y VGND VGND VPWR VPWR _14638_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16308_ _16320_/A _16320_/B VGND VGND VPWR VPWR _16308_/Y sky130_fd_sc_hd__nor2_1
X_14569_ _13009_/A _14568_/Y _13009_/A _14568_/Y VGND VGND VPWR VPWR _14571_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_118_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16239_ _16249_/B VGND VGND VPWR VPWR _16316_/A sky130_fd_sc_hd__buf_6
XFILLER_127_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08992_ _09518_/A _10134_/A _08752_/X _08868_/Y VGND VGND VPWR VPWR _08992_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09613_ _09613_/A _09613_/B VGND VGND VPWR VPWR _09613_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09544_ _09539_/A _09539_/B _09539_/X _09543_/X VGND VGND VPWR VPWR _09544_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09475_ _09450_/Y _09473_/X _09474_/X VGND VGND VPWR VPWR _09475_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08426_ _09213_/A VGND VGND VPWR VPWR _08714_/A sky130_fd_sc_hd__inv_2
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08357_ input26/X _08357_/B VGND VGND VPWR VPWR _08387_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08288_ input30/X _08341_/B _08342_/A _08344_/A VGND VGND VPWR VPWR _08339_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10250_ _10250_/A _10252_/B VGND VGND VPWR VPWR _10250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10181_ _10175_/Y _10179_/Y _10180_/Y VGND VGND VPWR VPWR _10182_/A sky130_fd_sc_hd__o21ai_1
XFILLER_94_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13940_ _14040_/A _13938_/X _13939_/X VGND VGND VPWR VPWR _13940_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15610_ _15539_/Y _15609_/A _15539_/A _15609_/Y _15595_/A VGND VGND VPWR VPWR _16040_/A
+ sky130_fd_sc_hd__a221o_1
X_13871_ _13871_/A _13872_/B VGND VGND VPWR VPWR _13873_/A sky130_fd_sc_hd__and2_1
XFILLER_74_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12822_ _12765_/X _12821_/Y _12765_/X _12821_/Y VGND VGND VPWR VPWR _12841_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15541_ _15536_/Y _15539_/Y _15540_/Y VGND VGND VPWR VPWR _15602_/A sky130_fd_sc_hd__o21ai_2
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _12711_/X _12752_/X _12711_/X _12752_/X VGND VGND VPWR VPWR _12768_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15472_ _12234_/Y _15471_/X _12234_/Y _15471_/X VGND VGND VPWR VPWR _15473_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11700_/X _11703_/X _11700_/X _11703_/X VGND VGND VPWR VPWR _11704_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_42_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _11776_/Y _14416_/X _11776_/Y _14416_/X VGND VGND VPWR VPWR _14424_/B sky130_fd_sc_hd__o2bb2a_1
X_12684_ _11328_/A _12675_/A _11328_/Y _12675_/Y VGND VGND VPWR VPWR _12685_/B sky130_fd_sc_hd__o22a_1
X_11635_ _11635_/A VGND VGND VPWR VPWR _11635_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14354_ _15881_/A _14250_/B _14250_/Y VGND VGND VPWR VPWR _14354_/Y sky130_fd_sc_hd__o21ai_1
X_11566_ _11468_/X _11565_/Y _11468_/X _11565_/Y VGND VGND VPWR VPWR _11567_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14285_ _14285_/A _15908_/A VGND VGND VPWR VPWR _14398_/B sky130_fd_sc_hd__or2_1
X_13305_ _13305_/A VGND VGND VPWR VPWR _13305_/Y sky130_fd_sc_hd__inv_2
X_10517_ _10517_/A VGND VGND VPWR VPWR _11794_/A sky130_fd_sc_hd__buf_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16024_ _15947_/Y _16023_/Y _15947_/Y _16023_/Y VGND VGND VPWR VPWR _16030_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13236_ _15066_/A VGND VGND VPWR VPWR _14473_/A sky130_fd_sc_hd__inv_2
X_11497_ _09997_/B _11496_/X _09997_/B _11496_/X VGND VGND VPWR VPWR _11498_/B sky130_fd_sc_hd__o2bb2a_1
X_10448_ _10450_/A VGND VGND VPWR VPWR _10448_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13167_ _13108_/X _13166_/Y _13108_/X _13166_/Y VGND VGND VPWR VPWR _13190_/B sky130_fd_sc_hd__a2bb2o_1
X_10379_ _11808_/A _10452_/B VGND VGND VPWR VPWR _10379_/Y sky130_fd_sc_hd__nand2_1
X_12118_ _13909_/A _12149_/B VGND VGND VPWR VPWR _12215_/A sky130_fd_sc_hd__and2_1
X_13098_ _14504_/A _13010_/B _13010_/Y VGND VGND VPWR VPWR _13098_/Y sky130_fd_sc_hd__a21oi_1
X_12049_ _12049_/A _12049_/B VGND VGND VPWR VPWR _12049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15808_ _15755_/Y _16197_/A _15807_/Y VGND VGND VPWR VPWR _15808_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15739_ _14917_/X _15738_/X _14917_/X _15738_/X VGND VGND VPWR VPWR _15740_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09260_ _09259_/X _08894_/Y _09259_/X _08894_/Y VGND VGND VPWR VPWR _10242_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09191_ _09429_/A _09191_/B VGND VGND VPWR VPWR _11667_/B sky130_fd_sc_hd__and2_1
XFILLER_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08975_ _08901_/X _08973_/X _11380_/B VGND VGND VPWR VPWR _08975_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09527_ _09527_/A _09527_/B VGND VGND VPWR VPWR _09528_/A sky130_fd_sc_hd__or2_1
XFILLER_52_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09458_ _09458_/A _09458_/B VGND VGND VPWR VPWR _09458_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08409_ _08409_/A VGND VGND VPWR VPWR _08409_/Y sky130_fd_sc_hd__inv_2
X_09389_ _09343_/X _09388_/X _09343_/X _09388_/X VGND VGND VPWR VPWR _10420_/B sky130_fd_sc_hd__a2bb2o_4
X_11420_ _11251_/X _11419_/X _11251_/X _11419_/X VGND VGND VPWR VPWR _11422_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11351_ _13889_/A _11352_/B VGND VGND VPWR VPWR _11353_/A sky130_fd_sc_hd__and2_1
X_10302_ _10454_/A _11226_/A VGND VGND VPWR VPWR _10303_/A sky130_fd_sc_hd__or2_1
XFILLER_106_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14070_ _14956_/A _13988_/B _13988_/Y _13991_/X VGND VGND VPWR VPWR _14070_/X sky130_fd_sc_hd__o2bb2a_1
X_11282_ _09438_/X _11281_/X _09438_/X _11281_/X VGND VGND VPWR VPWR _11283_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13021_ _14484_/A _13021_/B VGND VGND VPWR VPWR _13021_/X sky130_fd_sc_hd__or2_1
X_10233_ _10235_/A _10235_/B VGND VGND VPWR VPWR _10234_/A sky130_fd_sc_hd__or2_1
XFILLER_3_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10164_ _10113_/A _10113_/B _10114_/A VGND VGND VPWR VPWR _10167_/A sky130_fd_sc_hd__a21bo_1
XFILLER_121_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14972_ _14933_/Y _14971_/Y _14961_/Y VGND VGND VPWR VPWR _14972_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10095_ _09954_/Y _10094_/A _09954_/A _10094_/Y VGND VGND VPWR VPWR _11239_/A sky130_fd_sc_hd__a22o_2
X_13923_ _13842_/X _13922_/Y _13842_/X _13922_/Y VGND VGND VPWR VPWR _13943_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13854_ _13808_/Y _13852_/X _13853_/Y VGND VGND VPWR VPWR _13854_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12805_ _12853_/A _12853_/B VGND VGND VPWR VPWR _12805_/Y sky130_fd_sc_hd__nor2_1
X_15524_ _15524_/A _15524_/B VGND VGND VPWR VPWR _15524_/Y sky130_fd_sc_hd__nand2_1
X_10997_ _12162_/A _11115_/B VGND VGND VPWR VPWR _10997_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13785_ _13785_/A _13785_/B VGND VGND VPWR VPWR _13867_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _12780_/A _12780_/B VGND VGND VPWR VPWR _12736_/Y sky130_fd_sc_hd__nor2_1
X_15455_ _15455_/A _15455_/B VGND VGND VPWR VPWR _15455_/X sky130_fd_sc_hd__and2_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12667_/A VGND VGND VPWR VPWR _12667_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14406_ _12652_/Y _14405_/X _12652_/Y _14405_/X VGND VGND VPWR VPWR _14406_/Y sky130_fd_sc_hd__a2bb2oi_1
X_15386_ _15402_/A _15402_/B VGND VGND VPWR VPWR _15462_/A sky130_fd_sc_hd__and2_1
X_11618_ _11618_/A VGND VGND VPWR VPWR _11619_/B sky130_fd_sc_hd__inv_2
X_14337_ _14337_/B1 _14336_/Y _14337_/B1 _14336_/Y VGND VGND VPWR VPWR _14383_/A sky130_fd_sc_hd__a2bb2o_1
X_12598_ _14906_/A _11424_/B _11424_/Y VGND VGND VPWR VPWR _12599_/A sky130_fd_sc_hd__a21oi_1
XFILLER_11_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11549_ _12955_/A _11646_/B VGND VGND VPWR VPWR _11549_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14268_ _15863_/A _14268_/B VGND VGND VPWR VPWR _14268_/Y sky130_fd_sc_hd__nand2_1
X_16007_ _16042_/A _16042_/B VGND VGND VPWR VPWR _16007_/Y sky130_fd_sc_hd__nor2_1
X_14199_ _14110_/Y _14198_/X _14110_/Y _14198_/X VGND VGND VPWR VPWR _14200_/B sky130_fd_sc_hd__a2bb2oi_1
X_13219_ _13203_/X _13218_/Y _13203_/X _13218_/Y VGND VGND VPWR VPWR _13303_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08760_ _10133_/A VGND VGND VPWR VPWR _08760_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08691_ _08881_/A _08689_/X _08881_/B VGND VGND VPWR VPWR _08691_/X sky130_fd_sc_hd__o21ba_1
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09312_ _09312_/A _09312_/B VGND VGND VPWR VPWR _09312_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09243_ _09467_/B _09857_/A _09212_/Y _09242_/X VGND VGND VPWR VPWR _09243_/X sky130_fd_sc_hd__o22a_1
X_09174_ _09757_/A VGND VGND VPWR VPWR _09431_/A sky130_fd_sc_hd__buf_1
XFILLER_119_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08958_ _09538_/A _08635_/A _08637_/A VGND VGND VPWR VPWR _08958_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08889_ _08888_/Y _08864_/X _08888_/Y _08864_/X VGND VGND VPWR VPWR _08978_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10920_ _11027_/A _10917_/X _10919_/X VGND VGND VPWR VPWR _10920_/X sky130_fd_sc_hd__o21a_1
XFILLER_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10851_ _09265_/A _10850_/A _09268_/A _10850_/Y _10929_/A VGND VGND VPWR VPWR _12063_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _13530_/X _13569_/Y _13530_/X _13569_/Y VGND VGND VPWR VPWR _13573_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10782_ _10933_/A _10782_/B VGND VGND VPWR VPWR _13058_/A sky130_fd_sc_hd__or2_2
X_12521_ _12636_/A _12636_/B VGND VGND VPWR VPWR _14177_/A sky130_fd_sc_hd__and2_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A _15240_/B VGND VGND VPWR VPWR _15240_/Y sky130_fd_sc_hd__nand2_1
X_12452_ _12451_/Y _12368_/X _12390_/Y VGND VGND VPWR VPWR _12452_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11403_ _08952_/A _08952_/B _08952_/Y VGND VGND VPWR VPWR _11403_/X sky130_fd_sc_hd__o21a_1
X_15171_ _15171_/A _15425_/B VGND VGND VPWR VPWR _15171_/Y sky130_fd_sc_hd__nand2_1
X_12383_ _12381_/X _12383_/B VGND VGND VPWR VPWR _12383_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_126_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14122_ _14122_/A _14059_/X VGND VGND VPWR VPWR _14122_/X sky130_fd_sc_hd__or2b_1
X_11334_ _11519_/A _12376_/A _11333_/Y VGND VGND VPWR VPWR _11334_/X sky130_fd_sc_hd__a21o_1
X_14053_ _15458_/A _14027_/B _14027_/X _14052_/X VGND VGND VPWR VPWR _14053_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11265_ _11265_/A VGND VGND VPWR VPWR _11265_/Y sky130_fd_sc_hd__inv_2
X_13004_ _13004_/A VGND VGND VPWR VPWR _14504_/A sky130_fd_sc_hd__buf_1
X_10216_ _10216_/A VGND VGND VPWR VPWR _10216_/X sky130_fd_sc_hd__buf_1
XFILLER_121_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11196_ _11091_/X _11195_/X _11091_/X _11195_/X VGND VGND VPWR VPWR _11197_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10147_ _10147_/A _10147_/B VGND VGND VPWR VPWR _10147_/Y sky130_fd_sc_hd__nor2_1
X_14955_ _14952_/Y _14954_/X _14952_/Y _14954_/X VGND VGND VPWR VPWR _14956_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10078_ _10052_/X _10076_/X _10679_/B VGND VGND VPWR VPWR _10078_/X sky130_fd_sc_hd__o21a_1
X_13906_ _14614_/A _13851_/B _13851_/Y VGND VGND VPWR VPWR _13906_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14886_ _15540_/A _14916_/B VGND VGND VPWR VPWR _14886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13837_ _13837_/A _13837_/B VGND VGND VPWR VPWR _13837_/Y sky130_fd_sc_hd__nand2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13768_ _13768_/A _13768_/B VGND VGND VPWR VPWR _13768_/X sky130_fd_sc_hd__or2_1
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15507_ _15473_/A _15473_/B _15473_/Y VGND VGND VPWR VPWR _15507_/Y sky130_fd_sc_hd__o21ai_1
X_12719_ _12687_/A _12687_/B _12687_/Y _12718_/X VGND VGND VPWR VPWR _12719_/X sky130_fd_sc_hd__o2bb2a_1
X_15438_ _15362_/X _15438_/B VGND VGND VPWR VPWR _15438_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13699_ _13729_/A _13697_/X _13698_/X VGND VGND VPWR VPWR _13699_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15369_ _15369_/A _15345_/X VGND VGND VPWR VPWR _15369_/X sky130_fd_sc_hd__or2b_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09930_ _09928_/A _09928_/B _09929_/Y VGND VGND VPWR VPWR _09931_/B sky130_fd_sc_hd__o21ai_1
XFILLER_125_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09861_ _09861_/A _09861_/B VGND VGND VPWR VPWR _09924_/A sky130_fd_sc_hd__or2_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08812_ _09217_/A _09455_/B _08715_/X VGND VGND VPWR VPWR _08813_/A sky130_fd_sc_hd__o21ai_1
X_09792_ _09792_/A VGND VGND VPWR VPWR _09793_/B sky130_fd_sc_hd__inv_2
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08743_ _10009_/A _09525_/A VGND VGND VPWR VPWR _08743_/X sky130_fd_sc_hd__or2_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08674_ _09029_/A VGND VGND VPWR VPWR _08674_/Y sky130_fd_sc_hd__inv_2
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09226_ _09801_/A VGND VGND VPWR VPWR _09690_/A sky130_fd_sc_hd__inv_2
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09157_ _08710_/Y _09054_/Y _08740_/X VGND VGND VPWR VPWR _09158_/A sky130_fd_sc_hd__o21ai_1
X_09088_ _09088_/A VGND VGND VPWR VPWR _09088_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11050_ _15081_/A VGND VGND VPWR VPWR _12141_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10001_ _09569_/A _09999_/B _10001_/B1 _10000_/Y VGND VGND VPWR VPWR _10001_/X sky130_fd_sc_hd__o22a_1
XFILLER_103_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14740_ _14740_/A _14740_/B VGND VGND VPWR VPWR _14740_/X sky130_fd_sc_hd__or2_1
XFILLER_45_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11952_ _12992_/A _11901_/B _11901_/Y VGND VGND VPWR VPWR _11952_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10903_ _12049_/A VGND VGND VPWR VPWR _13832_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11883_ _11840_/A _11840_/B _11840_/Y VGND VGND VPWR VPWR _11883_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14671_ _15044_/A _12170_/Y _12092_/Y _14594_/X VGND VGND VPWR VPWR _14671_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16410_ _16406_/Y _16409_/Y _16349_/X _16349_/X _16402_/X VGND VGND VPWR VPWR _16411_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_83_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13622_ _13601_/Y _13619_/X _13621_/Y VGND VGND VPWR VPWR _13623_/A sky130_fd_sc_hd__o21ai_1
X_10834_ _10813_/X _10833_/X _10813_/X _10833_/X VGND VGND VPWR VPWR _10955_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16341_ input1/X VGND VGND VPWR VPWR _16361_/A sky130_fd_sc_hd__inv_2
X_13553_ _15036_/A _13518_/B _13518_/Y VGND VGND VPWR VPWR _13553_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12504_ _12412_/A _12412_/B _12412_/Y _12503_/X VGND VGND VPWR VPWR _12640_/B sky130_fd_sc_hd__o211a_1
X_10765_ _15212_/A _12043_/A VGND VGND VPWR VPWR _13008_/A sky130_fd_sc_hd__or2_1
XFILLER_40_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16272_ _16272_/A VGND VGND VPWR VPWR _16338_/A sky130_fd_sc_hd__buf_6
X_13484_ _10448_/Y _11767_/A _10387_/Y _13483_/X VGND VGND VPWR VPWR _13484_/X sky130_fd_sc_hd__o22a_1
X_10696_ _10812_/A _12693_/A _10695_/Y VGND VGND VPWR VPWR _10696_/X sky130_fd_sc_hd__a21o_1
X_15223_ _15196_/A _15196_/B _15196_/Y _15222_/X VGND VGND VPWR VPWR _15223_/X sky130_fd_sc_hd__a2bb2o_1
X_12435_ _13494_/A _12435_/B VGND VGND VPWR VPWR _12435_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12366_ _12364_/Y _12365_/Y _12286_/Y VGND VGND VPWR VPWR _12366_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15154_ _15125_/A _15125_/B _15125_/Y _15153_/X VGND VGND VPWR VPWR _15154_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14105_ _14105_/A _14105_/B VGND VGND VPWR VPWR _14105_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11317_ _11316_/Y _11141_/X _11150_/Y VGND VGND VPWR VPWR _11317_/X sky130_fd_sc_hd__o21a_1
X_12297_ _12295_/X _12297_/B VGND VGND VPWR VPWR _12297_/Y sky130_fd_sc_hd__nand2b_1
X_15085_ _10426_/A _12834_/Y _10422_/A _12831_/X VGND VGND VPWR VPWR _15087_/B sky130_fd_sc_hd__a22o_1
XFILLER_4_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14036_ _15400_/A _13941_/B _13941_/Y VGND VGND VPWR VPWR _14036_/X sky130_fd_sc_hd__o21a_1
X_11248_ _11248_/A _11074_/X VGND VGND VPWR VPWR _11248_/X sky130_fd_sc_hd__or2b_1
XFILLER_121_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11179_ _14061_/A _11179_/B VGND VGND VPWR VPWR _11179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15987_ _15854_/Y _15986_/X _15854_/Y _15986_/X VGND VGND VPWR VPWR _15987_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14938_ _15167_/A _14938_/B VGND VGND VPWR VPWR _14938_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14869_ _14778_/A _14778_/B _14778_/A _14778_/B VGND VGND VPWR VPWR _14869_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08390_ _08388_/Y _08389_/A _08388_/A _08389_/Y _08303_/A VGND VGND VPWR VPWR _09006_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09011_ _08904_/X _09023_/S _08604_/Y VGND VGND VPWR VPWR _09011_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09913_ _09913_/A _09913_/B VGND VGND VPWR VPWR _10949_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09844_ _09844_/A VGND VGND VPWR VPWR _09844_/Y sky130_fd_sc_hd__inv_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09775_ _09776_/A _09776_/B VGND VGND VPWR VPWR _09775_/Y sky130_fd_sc_hd__nor2_1
X_08726_ _08717_/A _08717_/B _08717_/X _08725_/Y VGND VGND VPWR VPWR _08726_/X sky130_fd_sc_hd__a22o_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08657_ _08657_/A VGND VGND VPWR VPWR _08657_/Y sky130_fd_sc_hd__inv_2
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08588_ _08587_/A _08343_/Y _08587_/Y _08343_/A VGND VGND VPWR VPWR _08589_/B sky130_fd_sc_hd__o22a_1
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10550_ _09700_/A _10549_/Y _09700_/Y _10549_/A _10959_/A VGND VGND VPWR VPWR _11853_/A
+ sky130_fd_sc_hd__o221a_1
X_10481_ _13628_/A _10533_/B VGND VGND VPWR VPWR _10481_/Y sky130_fd_sc_hd__nor2_1
X_09209_ _09209_/A _09209_/B VGND VGND VPWR VPWR _09857_/A sky130_fd_sc_hd__or2_2
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12220_ _12220_/A _12220_/B VGND VGND VPWR VPWR _12220_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12151_ _13905_/A _12151_/B VGND VGND VPWR VPWR _12151_/X sky130_fd_sc_hd__or2_1
XFILLER_123_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11102_ _12857_/A VGND VGND VPWR VPWR _15057_/A sky130_fd_sc_hd__clkbuf_2
X_12082_ _12082_/A _12082_/B VGND VGND VPWR VPWR _12082_/X sky130_fd_sc_hd__or2_1
X_15910_ _15910_/A VGND VGND VPWR VPWR _15978_/A sky130_fd_sc_hd__inv_2
X_11033_ _10870_/A _10870_/B _10870_/A _10870_/B VGND VGND VPWR VPWR _11033_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15841_ _14231_/A _15840_/Y _12618_/X VGND VGND VPWR VPWR _15841_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15772_ _14904_/A _14904_/B _14904_/Y VGND VGND VPWR VPWR _15773_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12984_ _13694_/A VGND VGND VPWR VPWR _14484_/A sky130_fd_sc_hd__inv_2
X_14723_ _15398_/A _14717_/B _14717_/X _14722_/X VGND VGND VPWR VPWR _14723_/X sky130_fd_sc_hd__o22a_1
X_11935_ _11915_/X _11934_/X _11915_/X _11934_/X VGND VGND VPWR VPWR _11983_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14654_ _14625_/Y _14652_/X _14653_/Y VGND VGND VPWR VPWR _14654_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13605_ _13605_/A _13605_/B VGND VGND VPWR VPWR _13605_/Y sky130_fd_sc_hd__nor2_1
X_11866_ _12774_/A _11917_/A _11865_/Y VGND VGND VPWR VPWR _11866_/Y sky130_fd_sc_hd__a21oi_1
X_14585_ _14585_/A _14585_/B VGND VGND VPWR VPWR _14585_/Y sky130_fd_sc_hd__nand2_1
X_11797_ _14428_/A _11790_/B _11790_/Y _11796_/X VGND VGND VPWR VPWR _11797_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10817_ _10078_/X _10816_/X _10078_/X _10816_/X VGND VGND VPWR VPWR _10818_/B sky130_fd_sc_hd__a2bb2o_1
X_16324_ _16324_/A _16324_/B VGND VGND VPWR VPWR _16324_/Y sky130_fd_sc_hd__nand2_1
X_10748_ _10633_/A _10747_/Y _10633_/A _10747_/Y VGND VGND VPWR VPWR _10749_/B sky130_fd_sc_hd__a2bb2o_1
X_13536_ _15038_/A _13515_/B _13515_/Y _13535_/X VGND VGND VPWR VPWR _13536_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16255_ _16255_/A _16255_/B VGND VGND VPWR VPWR _16255_/Y sky130_fd_sc_hd__nand2_1
X_13467_ _15289_/A _13139_/B _13139_/Y _13207_/X VGND VGND VPWR VPWR _13467_/X sky130_fd_sc_hd__o2bb2a_1
X_15206_ _15140_/A _15140_/B _15140_/Y VGND VGND VPWR VPWR _15206_/Y sky130_fd_sc_hd__o21ai_1
X_12418_ _12680_/A _12429_/B _15560_/A VGND VGND VPWR VPWR _12422_/A sky130_fd_sc_hd__o21ai_2
X_10679_ _10052_/X _10679_/B VGND VGND VPWR VPWR _10679_/X sky130_fd_sc_hd__and2b_1
X_16186_ _16262_/A _16328_/A VGND VGND VPWR VPWR _16186_/Y sky130_fd_sc_hd__nor2_1
X_13398_ _14092_/A VGND VGND VPWR VPWR _14095_/A sky130_fd_sc_hd__buf_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12349_ _14023_/A _12217_/B _12217_/Y VGND VGND VPWR VPWR _12349_/Y sky130_fd_sc_hd__o21ai_1
X_15137_ _15137_/A _15137_/B VGND VGND VPWR VPWR _15137_/Y sky130_fd_sc_hd__nand2_1
X_15068_ _15037_/X _15067_/X _15037_/X _15067_/X VGND VGND VPWR VPWR _15069_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14019_ _13950_/X _14018_/Y _13950_/X _14018_/Y VGND VGND VPWR VPWR _14055_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09560_ _08694_/A _09152_/A _09526_/Y _09559_/X VGND VGND VPWR VPWR _09560_/X sky130_fd_sc_hd__o22a_1
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09491_ _08798_/X _09468_/X _08798_/X _09468_/X VGND VGND VPWR VPWR _09492_/B sky130_fd_sc_hd__o2bb2a_1
X_08511_ _08567_/B VGND VGND VPWR VPWR _09791_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08442_ _08440_/A _08323_/Y _08440_/Y _08323_/A _08441_/X VGND VGND VPWR VPWR _08554_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08373_ input17/X _08254_/B _08327_/B _08372_/X VGND VGND VPWR VPWR _08440_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ _09808_/A _09503_/B _09817_/A _09817_/B _09826_/X VGND VGND VPWR VPWR _09827_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_19_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09758_ _09739_/A _09739_/B _09742_/A VGND VGND VPWR VPWR _10043_/A sky130_fd_sc_hd__a21bo_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08709_ _09330_/A _09476_/B VGND VGND VPWR VPWR _08709_/Y sky130_fd_sc_hd__nor2_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11791_/A _11720_/B VGND VGND VPWR VPWR _11720_/Y sky130_fd_sc_hd__nor2_1
X_09689_ _09689_/A _09689_/B VGND VGND VPWR VPWR _09692_/A sky130_fd_sc_hd__or2_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11649_/X _11651_/B VGND VGND VPWR VPWR _11651_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_30_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14370_ _15838_/A VGND VGND VPWR VPWR _14370_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10602_ _11882_/A _10639_/B VGND VGND VPWR VPWR _10602_/Y sky130_fd_sc_hd__nor2_1
X_11582_ _11632_/A VGND VGND VPWR VPWR _12789_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13321_ _13296_/A _13320_/Y _13296_/A _13320_/Y VGND VGND VPWR VPWR _13366_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10533_ _11846_/A _10533_/B VGND VGND VPWR VPWR _10533_/Y sky130_fd_sc_hd__nand2_1
X_16040_ _16040_/A _16040_/B VGND VGND VPWR VPWR _16040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13252_ _14422_/A VGND VGND VPWR VPWR _14728_/A sky130_fd_sc_hd__buf_1
X_10464_ _11857_/A _10556_/B VGND VGND VPWR VPWR _10464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13183_ _15329_/A _13182_/B _12045_/Y _13182_/Y VGND VGND VPWR VPWR _13183_/X sky130_fd_sc_hd__o2bb2a_1
X_12203_ _12201_/X _12203_/B VGND VGND VPWR VPWR _12203_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10395_ _09285_/Y _10394_/A _09285_/A _10394_/Y _09391_/A VGND VGND VPWR VPWR _10396_/A
+ sky130_fd_sc_hd__o221a_1
X_12134_ _12049_/A _12049_/B _12049_/Y VGND VGND VPWR VPWR _12134_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12065_ _12065_/A _12065_/B VGND VGND VPWR VPWR _12065_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11016_ _11016_/A VGND VGND VPWR VPWR _13547_/A sky130_fd_sc_hd__buf_1
X_15824_ _15706_/X _15822_/X _15834_/B VGND VGND VPWR VPWR _15824_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15755_ _16106_/A _15807_/B VGND VGND VPWR VPWR _15755_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12967_ _14668_/A _13031_/B VGND VGND VPWR VPWR _13050_/A sky130_fd_sc_hd__and2_1
XFILLER_18_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15686_ _15585_/Y _15684_/X _15685_/Y VGND VGND VPWR VPWR _15694_/A sky130_fd_sc_hd__o21a_1
X_14706_ _14650_/X _14705_/Y _14650_/X _14705_/Y VGND VGND VPWR VPWR _14728_/B sky130_fd_sc_hd__a2bb2o_1
X_12898_ _12845_/A _12845_/B _12845_/Y VGND VGND VPWR VPWR _12898_/Y sky130_fd_sc_hd__o21ai_1
X_11918_ _11916_/A _11916_/B _11916_/X _11917_/Y VGND VGND VPWR VPWR _11987_/B sky130_fd_sc_hd__a22o_1
X_14637_ _15333_/A _14647_/B VGND VGND VPWR VPWR _14637_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11849_ _13555_/A _11848_/B _11848_/X _11800_/X VGND VGND VPWR VPWR _11849_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _15216_/A _14507_/B _14507_/Y VGND VGND VPWR VPWR _14568_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16307_ _16252_/X _16306_/Y _16252_/X _16306_/Y VGND VGND VPWR VPWR _16320_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14499_ _15208_/A _14511_/B VGND VGND VPWR VPWR _14560_/A sky130_fd_sc_hd__and2_1
X_13519_ _13521_/A VGND VGND VPWR VPWR _15034_/A sky130_fd_sc_hd__buf_1
X_16238_ _16238_/A _16238_/B VGND VGND VPWR VPWR _16249_/B sky130_fd_sc_hd__or2_1
X_16169_ _16266_/B VGND VGND VPWR VPWR _16332_/A sky130_fd_sc_hd__buf_6
XFILLER_88_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08991_ _09478_/A VGND VGND VPWR VPWR _09518_/A sky130_fd_sc_hd__buf_1
XFILLER_96_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09612_ _09977_/A VGND VGND VPWR VPWR _09978_/A sky130_fd_sc_hd__buf_1
X_09543_ _09540_/A _09540_/B _09540_/X _09628_/B VGND VGND VPWR VPWR _09543_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09474_ _10010_/A _09474_/B VGND VGND VPWR VPWR _09474_/X sky130_fd_sc_hd__or2_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08425_ _08424_/A _08338_/Y _08424_/Y _08338_/A _08441_/A VGND VGND VPWR VPWR _09213_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08356_ _08354_/Y _08355_/A _08354_/A _08355_/Y _08303_/A VGND VGND VPWR VPWR _09225_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08287_ input29/X _08346_/B _08347_/A _08349_/A VGND VGND VPWR VPWR _08344_/A sky130_fd_sc_hd__o22a_1
XFILLER_20_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10180_ _10180_/A _10180_/B VGND VGND VPWR VPWR _10180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13870_ _13541_/X _13869_/Y _13541_/X _13869_/Y VGND VGND VPWR VPWR _13872_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12821_ _12766_/A _12766_/B _12766_/Y VGND VGND VPWR VPWR _12821_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15540_ _15540_/A _15540_/B VGND VGND VPWR VPWR _15540_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12752_ _12701_/A _12701_/B _12701_/Y VGND VGND VPWR VPWR _12752_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15471_ _15471_/A _15395_/X VGND VGND VPWR VPWR _15471_/X sky130_fd_sc_hd__or2b_1
XFILLER_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _15556_/A _11644_/B _11644_/X _11647_/Y VGND VGND VPWR VPWR _11703_/X sky130_fd_sc_hd__a22o_1
X_12683_ _12683_/A _12683_/B VGND VGND VPWR VPWR _12683_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14422_/A _14422_/B VGND VGND VPWR VPWR _14422_/Y sky130_fd_sc_hd__nor2_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _12442_/A _11634_/B VGND VGND VPWR VPWR _11634_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14353_ _14379_/A _15950_/A VGND VGND VPWR VPWR _14353_/X sky130_fd_sc_hd__and2_1
X_11565_ _14065_/A _11564_/B _11564_/Y VGND VGND VPWR VPWR _11565_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14284_ _12637_/X _14283_/X _12637_/X _14283_/X VGND VGND VPWR VPWR _14284_/X sky130_fd_sc_hd__a2bb2o_1
X_13304_ _13220_/Y _13302_/Y _13303_/Y VGND VGND VPWR VPWR _13305_/A sky130_fd_sc_hd__o21ai_2
X_10516_ _11836_/A VGND VGND VPWR VPWR _13609_/A sky130_fd_sc_hd__buf_1
X_11496_ _11496_/A _09788_/X VGND VGND VPWR VPWR _11496_/X sky130_fd_sc_hd__or2b_1
X_16023_ _15945_/X _16023_/B VGND VGND VPWR VPWR _16023_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_115_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13235_ _14736_/A _13294_/B VGND VGND VPWR VPWR _13235_/Y sky130_fd_sc_hd__nor2_1
X_10447_ _11804_/A VGND VGND VPWR VPWR _13518_/A sky130_fd_sc_hd__buf_1
XFILLER_123_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13166_ _15258_/A _13109_/B _13109_/Y VGND VGND VPWR VPWR _13166_/Y sky130_fd_sc_hd__o21ai_1
X_10378_ _10377_/A _10376_/Y _10377_/Y _10376_/A _10462_/A VGND VGND VPWR VPWR _10452_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13097_ _13101_/A VGND VGND VPWR VPWR _14567_/A sky130_fd_sc_hd__buf_1
X_12117_ _12060_/X _12116_/Y _12060_/X _12116_/Y VGND VGND VPWR VPWR _12149_/B sky130_fd_sc_hd__a2bb2o_1
X_12048_ _13832_/A _12049_/B VGND VGND VPWR VPWR _12048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15807_ _16106_/A _15807_/B VGND VGND VPWR VPWR _15807_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13999_ _13983_/X _13986_/X _13985_/B VGND VGND VPWR VPWR _13999_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15738_ _15542_/A _14918_/B _14918_/Y VGND VGND VPWR VPWR _15738_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15669_ _15669_/A _15669_/B VGND VGND VPWR VPWR _15669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09190_ _11667_/A _09190_/B VGND VGND VPWR VPWR _09190_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08974_ _08974_/A _08974_/B VGND VGND VPWR VPWR _11380_/B sky130_fd_sc_hd__or2_1
XFILLER_130_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09526_ _09526_/A VGND VGND VPWR VPWR _09526_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09457_ _09498_/A _09457_/B VGND VGND VPWR VPWR _09457_/Y sky130_fd_sc_hd__nor2_1
X_08408_ _09228_/A _08386_/Y _08407_/Y VGND VGND VPWR VPWR _08408_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09388_ _09359_/X _09387_/Y _09359_/X _09387_/Y VGND VGND VPWR VPWR _09388_/X sky130_fd_sc_hd__a2bb2o_1
X_08339_ _08339_/A VGND VGND VPWR VPWR _08339_/Y sky130_fd_sc_hd__inv_2
X_11350_ _11280_/X _11349_/X _11280_/X _11349_/X VGND VGND VPWR VPWR _11352_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10301_ _09112_/A _10300_/X _09112_/A _10300_/X VGND VGND VPWR VPWR _11226_/A sky130_fd_sc_hd__a2bb2o_2
X_13020_ _13080_/A _13018_/X _13019_/X VGND VGND VPWR VPWR _13020_/X sky130_fd_sc_hd__o21a_1
X_11281_ _09785_/A _09373_/A _09431_/X VGND VGND VPWR VPWR _11281_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10232_ _09297_/A _10230_/B _10231_/Y _10108_/Y VGND VGND VPWR VPWR _10235_/B sky130_fd_sc_hd__o22a_1
XFILLER_4_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10163_ _10163_/A _10163_/B VGND VGND VPWR VPWR _10163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14971_ _14971_/A _14971_/B VGND VGND VPWR VPWR _14971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10094_ _10094_/A VGND VGND VPWR VPWR _10094_/Y sky130_fd_sc_hd__inv_2
X_13922_ _14630_/A _13843_/B _13843_/Y VGND VGND VPWR VPWR _13922_/Y sky130_fd_sc_hd__o21ai_1
X_13853_ _14610_/A _13853_/B VGND VGND VPWR VPWR _13853_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12804_ _12777_/X _12803_/Y _12777_/X _12803_/Y VGND VGND VPWR VPWR _12853_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15523_ _15476_/X _15522_/Y _15476_/X _15522_/Y VGND VGND VPWR VPWR _15632_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10996_ _10947_/X _10995_/Y _10947_/X _10995_/Y VGND VGND VPWR VPWR _11115_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13784_ _13540_/X _13783_/Y _13540_/X _13783_/Y VGND VGND VPWR VPWR _13785_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12735_ _12717_/X _12734_/X _12717_/X _12734_/X VGND VGND VPWR VPWR _12780_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15454_ _15407_/X _15453_/X _15407_/X _15453_/X VGND VGND VPWR VPWR _15455_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _10677_/Y _12665_/Y _10566_/Y VGND VGND VPWR VPWR _12667_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14405_ _14290_/Y _14403_/X _14404_/Y VGND VGND VPWR VPWR _14405_/X sky130_fd_sc_hd__o21a_1
X_12597_ _14901_/A VGND VGND VPWR VPWR _14906_/A sky130_fd_sc_hd__buf_1
X_15385_ _15334_/X _15384_/X _15334_/X _15384_/X VGND VGND VPWR VPWR _15402_/B sky130_fd_sc_hd__a2bb2o_1
X_11617_ _11614_/X _11692_/A _11614_/A _11692_/A VGND VGND VPWR VPWR _11618_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14336_ _15872_/A _14259_/B _14259_/Y VGND VGND VPWR VPWR _14336_/Y sky130_fd_sc_hd__o21ai_1
X_11548_ _11501_/X _11547_/Y _11501_/X _11547_/Y VGND VGND VPWR VPWR _11646_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14267_ _14267_/A VGND VGND VPWR VPWR _14267_/Y sky130_fd_sc_hd__inv_2
X_11479_ _13872_/A VGND VGND VPWR VPWR _15107_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16006_ _15959_/X _16005_/Y _15959_/X _16005_/Y VGND VGND VPWR VPWR _16042_/B sky130_fd_sc_hd__a2bb2o_1
X_14198_ _14111_/A _14111_/B _14111_/Y VGND VGND VPWR VPWR _14198_/X sky130_fd_sc_hd__o21a_1
X_13218_ _13204_/A _13204_/B _13204_/Y VGND VGND VPWR VPWR _13218_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13149_ _13120_/X _13148_/Y _13120_/X _13148_/Y VGND VGND VPWR VPWR _13202_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08690_ _08690_/A _10118_/B VGND VGND VPWR VPWR _08881_/B sky130_fd_sc_hd__and2_1
XFILLER_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09311_ _09312_/A _09312_/B VGND VGND VPWR VPWR _09311_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09242_ _08597_/A _09856_/A _09216_/Y _09241_/X VGND VGND VPWR VPWR _09242_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09173_ _10010_/B _09165_/B _09166_/B VGND VGND VPWR VPWR _09757_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08957_ _08960_/A _08960_/B VGND VGND VPWR VPWR _08957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08888_ _09470_/A _08786_/B _08786_/Y VGND VGND VPWR VPWR _08888_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10850_ _10850_/A VGND VGND VPWR VPWR _10850_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09509_ _09498_/A _09498_/B _09498_/Y _09508_/X VGND VGND VPWR VPWR _09509_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10781_ _09657_/X _10780_/X _09657_/X _10780_/X VGND VGND VPWR VPWR _10782_/B sky130_fd_sc_hd__a2bb2oi_1
X_12520_ _12519_/A _12519_/B _12519_/Y _12503_/X VGND VGND VPWR VPWR _12636_/B sky130_fd_sc_hd__o211a_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _13974_/A _12451_/B VGND VGND VPWR VPWR _12451_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15170_ _15168_/X _15169_/Y _15168_/X _15169_/Y VGND VGND VPWR VPWR _15425_/B sky130_fd_sc_hd__a2bb2o_1
X_11402_ _11399_/Y _11401_/Y _11399_/A _11401_/A _12606_/B VGND VGND VPWR VPWR _13397_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_126_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14121_ _14115_/X _14118_/Y _14876_/A _14120_/Y VGND VGND VPWR VPWR _14121_/X sky130_fd_sc_hd__o22a_1
X_12382_ _12382_/A _12382_/B VGND VGND VPWR VPWR _12383_/B sky130_fd_sc_hd__or2_1
XFILLER_125_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11333_ _11519_/A _12376_/A VGND VGND VPWR VPWR _11333_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14052_ _15461_/A _14031_/B _14031_/X _14051_/X VGND VGND VPWR VPWR _14052_/X sky130_fd_sc_hd__o22a_1
XFILLER_4_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11264_ _09431_/A _09180_/B _09180_/Y VGND VGND VPWR VPWR _11265_/A sky130_fd_sc_hd__o21ai_1
XFILLER_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13003_ _13676_/A _13012_/B VGND VGND VPWR VPWR _13003_/Y sky130_fd_sc_hd__nor2_1
X_10215_ _10215_/A VGND VGND VPWR VPWR _10454_/A sky130_fd_sc_hd__buf_6
X_11195_ _11195_/A _11092_/X VGND VGND VPWR VPWR _11195_/X sky130_fd_sc_hd__or2b_1
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10146_ _10131_/A _10131_/B _10132_/B VGND VGND VPWR VPWR _10147_/B sky130_fd_sc_hd__a21bo_1
X_14954_ _14834_/X _14953_/Y _14851_/Y VGND VGND VPWR VPWR _14954_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10077_ _10077_/A _10077_/B VGND VGND VPWR VPWR _10679_/B sky130_fd_sc_hd__or2_1
X_13905_ _13905_/A VGND VGND VPWR VPWR _15410_/A sky130_fd_sc_hd__buf_1
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14885_ _14821_/X _14884_/X _14821_/X _14884_/X VGND VGND VPWR VPWR _14916_/B sky130_fd_sc_hd__a2bb2o_1
X_13836_ _14643_/A _13837_/B VGND VGND VPWR VPWR _13836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13767_ _13812_/A _13765_/X _13766_/X VGND VGND VPWR VPWR _13767_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10979_ _12176_/A _11140_/B _10978_/Y VGND VGND VPWR VPWR _10980_/A sky130_fd_sc_hd__o21ai_2
XFILLER_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15506_ _15542_/A _15542_/B VGND VGND VPWR VPWR _15600_/A sky130_fd_sc_hd__and2_1
X_12718_ _12689_/A _12689_/B _12689_/Y _12717_/X VGND VGND VPWR VPWR _12718_/X sky130_fd_sc_hd__o2bb2a_1
X_15437_ _15437_/A _15437_/B VGND VGND VPWR VPWR _15437_/X sky130_fd_sc_hd__and2_1
X_13698_ _13698_/A _13698_/B VGND VGND VPWR VPWR _13698_/X sky130_fd_sc_hd__or2_1
XFILLER_31_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12649_ _12649_/A _12649_/B VGND VGND VPWR VPWR _12651_/B sky130_fd_sc_hd__or2_1
XFILLER_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15368_ _15414_/A _15414_/B VGND VGND VPWR VPWR _15444_/A sky130_fd_sc_hd__and2_1
XFILLER_116_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14319_ _13436_/X _14318_/X _13436_/X _14318_/X VGND VGND VPWR VPWR _14320_/B sky130_fd_sc_hd__a2bb2oi_1
X_15299_ _15349_/A _15349_/B VGND VGND VPWR VPWR _15363_/A sky130_fd_sc_hd__and2_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09860_ _09860_/A _09914_/A VGND VGND VPWR VPWR _09861_/B sky130_fd_sc_hd__or2_1
XFILLER_98_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08811_ _09456_/A VGND VGND VPWR VPWR _09496_/A sky130_fd_sc_hd__buf_1
X_09791_ _09791_/A _09791_/B _09791_/C VGND VGND VPWR VPWR _09792_/A sky130_fd_sc_hd__or3_2
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08742_ _08742_/A VGND VGND VPWR VPWR _08742_/Y sky130_fd_sc_hd__inv_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08673_ _10228_/A _10098_/A VGND VGND VPWR VPWR _09029_/A sky130_fd_sc_hd__or2_1
XFILLER_93_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09225_ _09225_/A _09225_/B VGND VGND VPWR VPWR _09801_/A sky130_fd_sc_hd__or2_1
XFILLER_21_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09156_ _09525_/B _09156_/B VGND VGND VPWR VPWR _09156_/X sky130_fd_sc_hd__or2_1
X_09087_ _09551_/B _09034_/B _09035_/B VGND VGND VPWR VPWR _09088_/A sky130_fd_sc_hd__a21bo_1
XFILLER_107_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10000_ _10000_/A VGND VGND VPWR VPWR _10000_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09989_ _09989_/A _09990_/B VGND VGND VPWR VPWR _09989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11951_ _13078_/A _11972_/B VGND VGND VPWR VPWR _11951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10902_ _10907_/A _10902_/B VGND VGND VPWR VPWR _12049_/A sky130_fd_sc_hd__nand2b_1
XFILLER_84_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11882_ _11882_/A _11901_/B VGND VGND VPWR VPWR _11882_/Y sky130_fd_sc_hd__nor2_1
X_14670_ _14596_/A _14596_/B _14593_/X _14596_/Y VGND VGND VPWR VPWR _14670_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13621_ _15137_/A _13621_/B VGND VGND VPWR VPWR _13621_/Y sky130_fd_sc_hd__nand2_1
X_10833_ _10964_/A _12691_/A _10832_/Y VGND VGND VPWR VPWR _10833_/X sky130_fd_sc_hd__a21o_1
X_16340_ _16278_/Y _16339_/X _16278_/Y _16339_/X VGND VGND VPWR VPWR _16392_/A sky130_fd_sc_hd__a2bb2o_1
X_10764_ _13753_/A VGND VGND VPWR VPWR _11063_/A sky130_fd_sc_hd__inv_2
X_13552_ _13552_/A VGND VGND VPWR VPWR _13552_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12503_ _12503_/A VGND VGND VPWR VPWR _12503_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16271_ _16154_/Y _16269_/X _16270_/Y VGND VGND VPWR VPWR _16271_/X sky130_fd_sc_hd__o21a_1
X_13483_ _10365_/Y _11753_/A _10316_/Y _13482_/X VGND VGND VPWR VPWR _13483_/X sky130_fd_sc_hd__o22a_1
X_10695_ _10812_/A _11992_/A VGND VGND VPWR VPWR _10695_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15222_ _15199_/A _15199_/B _15199_/Y _15221_/X VGND VGND VPWR VPWR _15222_/X sky130_fd_sc_hd__a2bb2o_1
X_12434_ _13457_/A _12424_/Y _12432_/A _12431_/X _12433_/X VGND VGND VPWR VPWR _12434_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_126_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12365_ _12365_/A VGND VGND VPWR VPWR _12365_/Y sky130_fd_sc_hd__inv_2
X_15153_ _15128_/A _15128_/B _15128_/Y _15152_/X VGND VGND VPWR VPWR _15153_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14104_ _14052_/X _14103_/X _14052_/X _14103_/X VGND VGND VPWR VPWR _14104_/Y sky130_fd_sc_hd__a2bb2oi_1
X_15084_ _15084_/A _15084_/B VGND VGND VPWR VPWR _15084_/Y sky130_fd_sc_hd__nand2_1
X_11316_ _12270_/A _11316_/B VGND VGND VPWR VPWR _11316_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14035_ _14035_/A _14035_/B VGND VGND VPWR VPWR _14035_/X sky130_fd_sc_hd__and2_1
X_12296_ _13889_/A _12296_/B VGND VGND VPWR VPWR _12297_/B sky130_fd_sc_hd__or2_1
XFILLER_4_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11247_ _12234_/A _13935_/B VGND VGND VPWR VPWR _11247_/X sky130_fd_sc_hd__or2_1
XFILLER_122_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11178_ _11095_/X _11177_/X _11095_/X _11177_/X VGND VGND VPWR VPWR _11179_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10129_ _10129_/A _10129_/B VGND VGND VPWR VPWR _10130_/B sky130_fd_sc_hd__or2_1
X_15986_ _15983_/Y _15985_/X _15983_/Y _15985_/X VGND VGND VPWR VPWR _15986_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14937_ _12439_/A _14936_/X _12439_/A _14936_/X VGND VGND VPWR VPWR _14938_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14868_ _14868_/A VGND VGND VPWR VPWR _15548_/A sky130_fd_sc_hd__buf_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13819_ _13761_/X _13818_/X _13761_/X _13818_/X VGND VGND VPWR VPWR _13845_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14799_ _15461_/A VGND VGND VPWR VPWR _14802_/A sky130_fd_sc_hd__buf_1
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16469_ _08229_/A _16469_/D VGND VGND VPWR VPWR _16469_/Q sky130_fd_sc_hd__dfxtp_1
X_09010_ _09496_/A _09024_/S _09221_/B VGND VGND VPWR VPWR _09023_/S sky130_fd_sc_hd__a21oi_1
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09912_ _09913_/A _09913_/B VGND VGND VPWR VPWR _10949_/B sky130_fd_sc_hd__and2_1
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09843_ _09843_/A _09843_/B VGND VGND VPWR VPWR _10490_/B sky130_fd_sc_hd__nor2_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _10077_/A _09772_/Y _09773_/Y VGND VGND VPWR VPWR _09776_/B sky130_fd_sc_hd__o21ai_1
XFILLER_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08725_ _08718_/Y _08723_/X _08724_/X VGND VGND VPWR VPWR _08725_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08656_ _08656_/A _09684_/A VGND VGND VPWR VPWR _08657_/A sky130_fd_sc_hd__or2_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08587_ _08587_/A VGND VGND VPWR VPWR _08587_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_26_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09208_ _14061_/A VGND VGND VPWR VPWR _15443_/A sky130_fd_sc_hd__buf_1
X_10480_ _10435_/X _10479_/X _10435_/X _10479_/X VGND VGND VPWR VPWR _10533_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09139_ _09531_/B _09037_/B _09038_/B VGND VGND VPWR VPWR _09140_/A sky130_fd_sc_hd__a21bo_1
XFILLER_118_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12150_ _12215_/A _12148_/X _12149_/X VGND VGND VPWR VPWR _12150_/X sky130_fd_sc_hd__o21a_1
X_11101_ _13712_/A VGND VGND VPWR VPWR _12857_/A sky130_fd_sc_hd__buf_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12081_ _12169_/A VGND VGND VPWR VPWR _12780_/A sky130_fd_sc_hd__buf_1
XFILLER_1_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11032_ _15072_/A VGND VGND VPWR VPWR _13913_/A sky130_fd_sc_hd__buf_1
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15840_ _15840_/A VGND VGND VPWR VPWR _15840_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15771_ _16086_/A VGND VGND VPWR VPWR _16089_/A sky130_fd_sc_hd__clkbuf_2
X_12983_ _14480_/A _13023_/B VGND VGND VPWR VPWR _13070_/A sky130_fd_sc_hd__and2_1
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14722_ _13936_/X _14720_/Y _14721_/Y VGND VGND VPWR VPWR _14722_/X sky130_fd_sc_hd__o21a_1
X_11934_ _10666_/X _11985_/B _10666_/X _11985_/B VGND VGND VPWR VPWR _11934_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14653_ _15339_/A _14653_/B VGND VGND VPWR VPWR _14653_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13604_ _13574_/Y _13603_/Y _13574_/Y _13603_/Y VGND VGND VPWR VPWR _13605_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11865_ _12774_/A _11917_/A VGND VGND VPWR VPWR _11865_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14584_ _14546_/Y _14582_/X _14583_/Y VGND VGND VPWR VPWR _14584_/X sky130_fd_sc_hd__o21a_1
X_11796_ _12827_/A _11794_/B _11794_/X _11795_/X VGND VGND VPWR VPWR _11796_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10816_ _10049_/X _10816_/B VGND VGND VPWR VPWR _10816_/X sky130_fd_sc_hd__and2b_1
X_16323_ _16305_/Y _16321_/X _16322_/Y VGND VGND VPWR VPWR _16323_/X sky130_fd_sc_hd__o21a_1
X_10747_ _12997_/A _10635_/B _10635_/Y VGND VGND VPWR VPWR _10747_/Y sky130_fd_sc_hd__o21ai_1
X_13535_ _15036_/A _13518_/B _13518_/Y _13534_/X VGND VGND VPWR VPWR _13535_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16254_ _16221_/Y _16252_/X _16253_/Y VGND VGND VPWR VPWR _16254_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13466_ _12428_/A _12680_/B _12680_/Y _12721_/X VGND VGND VPWR VPWR _13466_/Y sky130_fd_sc_hd__o2bb2ai_1
X_10678_ _10677_/Y _10557_/X _10566_/Y VGND VGND VPWR VPWR _10678_/X sky130_fd_sc_hd__o21a_1
X_15205_ _15205_/A _15205_/B VGND VGND VPWR VPWR _15205_/Y sky130_fd_sc_hd__nand2_1
X_12417_ _12680_/A _12429_/B VGND VGND VPWR VPWR _15560_/A sky130_fd_sc_hd__nand2_1
X_16185_ _16262_/B VGND VGND VPWR VPWR _16328_/A sky130_fd_sc_hd__buf_6
X_13397_ _13397_/A VGND VGND VPWR VPWR _14092_/A sky130_fd_sc_hd__inv_2
XFILLER_114_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12348_ _12351_/A _12351_/B VGND VGND VPWR VPWR _12348_/Y sky130_fd_sc_hd__nor2_1
X_15136_ _15090_/X _15135_/Y _15090_/X _15135_/Y VGND VGND VPWR VPWR _15137_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12279_ _12784_/A _12372_/A _12278_/Y VGND VGND VPWR VPWR _12279_/Y sky130_fd_sc_hd__a21oi_1
X_15067_ _15067_/A _15038_/X VGND VGND VPWR VPWR _15067_/X sky130_fd_sc_hd__or2b_1
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14018_ _15410_/A _13951_/B _13951_/Y VGND VGND VPWR VPWR _14018_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15969_ _15966_/A _15966_/B _15966_/Y _15968_/X VGND VGND VPWR VPWR _15969_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09490_ _09490_/A _09490_/B VGND VGND VPWR VPWR _09490_/Y sky130_fd_sc_hd__nor2_1
X_08510_ _08656_/A VGND VGND VPWR VPWR _08567_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08441_ _08441_/A VGND VGND VPWR VPWR _08441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08372_ input16/X _08257_/B _08332_/B _08429_/A VGND VGND VPWR VPWR _08372_/X sky130_fd_sc_hd__o22a_1
XFILLER_23_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ _09826_/A _09826_/B VGND VGND VPWR VPWR _09826_/X sky130_fd_sc_hd__or2_1
X_09757_ _09757_/A VGND VGND VPWR VPWR _09785_/A sky130_fd_sc_hd__inv_2
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _09448_/A _08755_/A VGND VGND VPWR VPWR _08708_/Y sky130_fd_sc_hd__nor2_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _08632_/X _09690_/B _08632_/X _09690_/B VGND VGND VPWR VPWR _09689_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08660_/A _08639_/B VGND VGND VPWR VPWR _09459_/B sky130_fd_sc_hd__or2_2
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11650_ _12445_/A _11650_/B VGND VGND VPWR VPWR _11651_/B sky130_fd_sc_hd__or2_1
XFILLER_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10601_ _10528_/X _10600_/Y _10528_/X _10600_/Y VGND VGND VPWR VPWR _10639_/B sky130_fd_sc_hd__a2bb2o_1
X_11581_ _13133_/A VGND VGND VPWR VPWR _11632_/A sky130_fd_sc_hd__buf_1
X_13320_ _14738_/A _13297_/B _13297_/Y VGND VGND VPWR VPWR _13320_/Y sky130_fd_sc_hd__o21ai_1
X_10532_ _10488_/Y _10530_/X _10531_/Y VGND VGND VPWR VPWR _10532_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13251_ _15075_/A VGND VGND VPWR VPWR _14422_/A sky130_fd_sc_hd__inv_2
XFILLER_10_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10463_ _10461_/A _10460_/Y _10461_/Y _10460_/A _10976_/A VGND VGND VPWR VPWR _10556_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13182_ _13832_/A _13182_/B VGND VGND VPWR VPWR _13182_/Y sky130_fd_sc_hd__nor2_1
X_12202_ _13893_/A _12202_/B VGND VGND VPWR VPWR _12203_/B sky130_fd_sc_hd__or2_1
XFILLER_89_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10394_ _10394_/A VGND VGND VPWR VPWR _10394_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12133_ _12139_/A _12139_/B VGND VGND VPWR VPWR _12230_/A sky130_fd_sc_hd__and2_1
XFILLER_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12064_ _12020_/Y _12062_/X _12063_/Y VGND VGND VPWR VPWR _12064_/X sky130_fd_sc_hd__o21a_1
X_11015_ _13901_/A _11092_/B VGND VGND VPWR VPWR _11195_/A sky130_fd_sc_hd__and2_1
XFILLER_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15823_ _16125_/A _15823_/B VGND VGND VPWR VPWR _15834_/B sky130_fd_sc_hd__or2_1
XFILLER_65_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15754_ _15674_/X _15753_/Y _15674_/X _15753_/Y VGND VGND VPWR VPWR _15807_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14705_ _15337_/A _14651_/B _14651_/Y VGND VGND VPWR VPWR _14705_/Y sky130_fd_sc_hd__o21ai_1
X_12966_ _12943_/X _12965_/Y _12943_/X _12965_/Y VGND VGND VPWR VPWR _13031_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15685_ _15685_/A _15685_/B VGND VGND VPWR VPWR _15685_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12897_ _12932_/A VGND VGND VPWR VPWR _14464_/A sky130_fd_sc_hd__buf_1
X_11917_ _11917_/A VGND VGND VPWR VPWR _11917_/Y sky130_fd_sc_hd__inv_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14574_/X _14635_/Y _14574_/X _14635_/Y VGND VGND VPWR VPWR _14647_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11848_ _11848_/A _11848_/B VGND VGND VPWR VPWR _11848_/X sky130_fd_sc_hd__and2_1
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14567_ _14567_/A VGND VGND VPWR VPWR _15270_/A sky130_fd_sc_hd__buf_1
XFILLER_14_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16306_ _16253_/A _16320_/A _16253_/Y VGND VGND VPWR VPWR _16306_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11779_ _11779_/A VGND VGND VPWR VPWR _12766_/A sky130_fd_sc_hd__buf_1
X_13518_ _13518_/A _13518_/B VGND VGND VPWR VPWR _13518_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14498_ _14459_/X _14497_/Y _14459_/X _14497_/Y VGND VGND VPWR VPWR _14511_/B sky130_fd_sc_hd__a2bb2o_1
X_16237_ _15789_/Y _16236_/X _15789_/Y _16236_/X VGND VGND VPWR VPWR _16238_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_127_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13449_ _13449_/A _13449_/B VGND VGND VPWR VPWR _13449_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16168_ _16192_/A _16168_/B VGND VGND VPWR VPWR _16266_/B sky130_fd_sc_hd__or2_1
X_15119_ _15119_/A _15119_/B VGND VGND VPWR VPWR _15119_/Y sky130_fd_sc_hd__nand2_1
X_16099_ _16099_/A _16099_/B VGND VGND VPWR VPWR _16099_/Y sky130_fd_sc_hd__nand2_1
X_08990_ _09478_/B _08989_/Y _08514_/Y _08695_/Y VGND VGND VPWR VPWR _08990_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09611_ _09509_/X _09610_/X _09509_/X _09610_/X VGND VGND VPWR VPWR _09977_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09542_ _09629_/B VGND VGND VPWR VPWR _09628_/B sky130_fd_sc_hd__inv_2
XFILLER_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09473_ _09451_/Y _09471_/X _09472_/X VGND VGND VPWR VPWR _09473_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08424_ _08424_/A VGND VGND VPWR VPWR _08424_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08355_ _08355_/A VGND VGND VPWR VPWR _08355_/Y sky130_fd_sc_hd__inv_2
X_08286_ input28/X _08352_/B _08353_/A _08355_/A VGND VGND VPWR VPWR _08349_/A sky130_fd_sc_hd__o22a_1
XFILLER_20_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09809_ _08844_/A _09230_/A _09459_/Y _09826_/A VGND VGND VPWR VPWR _09809_/X sky130_fd_sc_hd__o22a_1
XFILLER_101_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12820_ _12843_/A _12843_/B VGND VGND VPWR VPWR _12820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12751_ _12770_/A _12770_/B VGND VGND VPWR VPWR _12751_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15470_ _15470_/A _15470_/B VGND VGND VPWR VPWR _15470_/Y sky130_fd_sc_hd__nand2_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _13978_/A VGND VGND VPWR VPWR _15556_/A sky130_fd_sc_hd__buf_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12682_ _11533_/A _12677_/A _11533_/Y _12677_/Y VGND VGND VPWR VPWR _12683_/B sky130_fd_sc_hd__o22a_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14421_ _11771_/Y _14417_/X _11771_/Y _14417_/X VGND VGND VPWR VPWR _14422_/B sky130_fd_sc_hd__o2bb2a_1
X_11633_ _11632_/A _11632_/B _11632_/Y VGND VGND VPWR VPWR _11633_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14352_ _14352_/A _14352_/B VGND VGND VPWR VPWR _15950_/A sky130_fd_sc_hd__or2_1
X_11564_ _14065_/A _11564_/B VGND VGND VPWR VPWR _11564_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14283_ _14283_/A _12638_/X VGND VGND VPWR VPWR _14283_/X sky130_fd_sc_hd__or2b_1
X_13303_ _14771_/A _13303_/B VGND VGND VPWR VPWR _13303_/Y sky130_fd_sc_hd__nand2_1
X_11495_ _11493_/Y _11494_/Y _11343_/Y VGND VGND VPWR VPWR _11495_/X sky130_fd_sc_hd__o21a_1
X_10515_ _09403_/X _08931_/Y _08931_/A _10514_/Y _11595_/A VGND VGND VPWR VPWR _11836_/A
+ sky130_fd_sc_hd__a221o_2
X_16022_ _16032_/A _16032_/B VGND VGND VPWR VPWR _16022_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13234_ _13197_/X _13233_/Y _13197_/X _13233_/Y VGND VGND VPWR VPWR _13294_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10446_ _09970_/A _10444_/Y _09970_/Y _10444_/A _10959_/A VGND VGND VPWR VPWR _11804_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13165_ _13192_/A _13192_/B VGND VGND VPWR VPWR _13165_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10377_ _10377_/A VGND VGND VPWR VPWR _10377_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13096_ _13096_/A VGND VGND VPWR VPWR _13096_/X sky130_fd_sc_hd__buf_1
X_12116_ _13194_/A _12061_/B _12061_/Y VGND VGND VPWR VPWR _12116_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12047_ _11064_/A _12046_/X _11064_/A _12046_/X VGND VGND VPWR VPWR _12049_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15806_ _15802_/Y _16207_/A _15805_/Y VGND VGND VPWR VPWR _16197_/A sky130_fd_sc_hd__o21ai_2
XFILLER_92_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13998_ _15425_/A _13971_/A _13972_/Y _13997_/Y VGND VGND VPWR VPWR _13998_/X sky130_fd_sc_hd__o22a_1
X_15737_ _16112_/A _15813_/B VGND VGND VPWR VPWR _15737_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12949_ _14944_/A _12949_/B VGND VGND VPWR VPWR _12949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15668_ _15654_/X _15666_/X _15788_/B VGND VGND VPWR VPWR _15668_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14619_ _14583_/A _14583_/B _14583_/Y VGND VGND VPWR VPWR _14619_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15599_ _15681_/A _15681_/B VGND VGND VPWR VPWR _15599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08973_ _08907_/X _08971_/X _11387_/B VGND VGND VPWR VPWR _08973_/X sky130_fd_sc_hd__o21a_1
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09525_ _09525_/A _09525_/B VGND VGND VPWR VPWR _09526_/A sky130_fd_sc_hd__or2_1
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09456_ _09456_/A _09456_/B VGND VGND VPWR VPWR _09456_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08407_ _09006_/A _08403_/Y _09459_/A VGND VGND VPWR VPWR _08407_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09387_ _09429_/B _11577_/A _09364_/X _11579_/A VGND VGND VPWR VPWR _09387_/Y sky130_fd_sc_hd__a22oi_1
X_08338_ _08338_/A VGND VGND VPWR VPWR _08338_/Y sky130_fd_sc_hd__inv_2
X_08269_ _08269_/A input12/X VGND VGND VPWR VPWR _08353_/A sky130_fd_sc_hd__nor2_1
X_11280_ _14663_/A _11279_/B _11279_/X _11104_/X VGND VGND VPWR VPWR _11280_/X sky130_fd_sc_hd__o22a_1
X_10300_ _09717_/A _09113_/B _09113_/Y VGND VGND VPWR VPWR _10300_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10231_ _10231_/A VGND VGND VPWR VPWR _10231_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10162_ _08810_/B _10127_/B _10128_/B VGND VGND VPWR VPWR _10163_/B sky130_fd_sc_hd__a21bo_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14970_ _14935_/X _14949_/A _14948_/X VGND VGND VPWR VPWR _14970_/Y sky130_fd_sc_hd__o21ai_1
X_10093_ _10055_/A _10055_/B _10055_/X VGND VGND VPWR VPWR _10094_/A sky130_fd_sc_hd__a21bo_1
XFILLER_120_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13921_ _13921_/A VGND VGND VPWR VPWR _15402_/A sky130_fd_sc_hd__buf_1
XFILLER_75_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13852_ _13811_/Y _13850_/X _13851_/Y VGND VGND VPWR VPWR _13852_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12803_ _12778_/A _12778_/B _12778_/Y VGND VGND VPWR VPWR _12803_/Y sky130_fd_sc_hd__o21ai_1
X_13783_ _15051_/A _13500_/B _13500_/Y VGND VGND VPWR VPWR _13783_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15522_ _15464_/A _15464_/B _15464_/Y VGND VGND VPWR VPWR _15522_/Y sky130_fd_sc_hd__o21ai_1
X_10995_ _13705_/A _11122_/B _10994_/Y VGND VGND VPWR VPWR _10995_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _12689_/A _12689_/B _12689_/Y VGND VGND VPWR VPWR _12734_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15453_ _15453_/A _15408_/X VGND VGND VPWR VPWR _15453_/X sky130_fd_sc_hd__or2b_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12665_/A VGND VGND VPWR VPWR _12665_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14404_ _15982_/A _14404_/B VGND VGND VPWR VPWR _14404_/Y sky130_fd_sc_hd__nand2_1
X_12596_ _14083_/A VGND VGND VPWR VPWR _14901_/A sky130_fd_sc_hd__buf_1
X_15384_ _15384_/A _15335_/X VGND VGND VPWR VPWR _15384_/X sky130_fd_sc_hd__or2b_1
X_11616_ _11615_/Y _11522_/X _11531_/X VGND VGND VPWR VPWR _11692_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14335_ _14385_/A _15956_/A VGND VGND VPWR VPWR _14335_/X sky130_fd_sc_hd__and2_1
X_11547_ _13974_/A _11641_/B _11546_/Y VGND VGND VPWR VPWR _11547_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16005_ _15927_/X _16005_/B VGND VGND VPWR VPWR _16005_/Y sky130_fd_sc_hd__nand2b_1
X_14266_ _14203_/Y _14264_/Y _14265_/Y VGND VGND VPWR VPWR _14267_/A sky130_fd_sc_hd__o21ai_2
XFILLER_109_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11478_ _12442_/A VGND VGND VPWR VPWR _13872_/A sky130_fd_sc_hd__buf_1
XFILLER_124_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14197_ _15863_/A _14268_/B VGND VGND VPWR VPWR _14197_/Y sky130_fd_sc_hd__nor2_1
X_13217_ _14754_/A VGND VGND VPWR VPWR _14771_/A sky130_fd_sc_hd__buf_1
X_10429_ _12827_/A _10429_/B VGND VGND VPWR VPWR _10429_/X sky130_fd_sc_hd__and2_1
XFILLER_111_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13148_ _15240_/A _13121_/B _13121_/Y VGND VGND VPWR VPWR _13148_/Y sky130_fd_sc_hd__o21ai_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13079_ _13762_/A VGND VGND VPWR VPWR _15258_/A sky130_fd_sc_hd__buf_1
XFILLER_66_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09310_ _09946_/A _09308_/Y _09309_/Y VGND VGND VPWR VPWR _09312_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09241_ _08610_/A _09803_/A _09220_/Y _09240_/X VGND VGND VPWR VPWR _09241_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09172_ _09754_/A VGND VGND VPWR VPWR _09430_/A sky130_fd_sc_hd__buf_1
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08956_ _08954_/Y _08955_/Y _08954_/Y _08955_/Y VGND VGND VPWR VPWR _08960_/B sky130_fd_sc_hd__o2bb2a_1
X_08887_ _08687_/X _08886_/Y _08687_/X _08886_/Y VGND VGND VPWR VPWR _08978_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09508_ _09500_/A _09500_/B _09500_/Y _09507_/X VGND VGND VPWR VPWR _09508_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10780_ _09987_/A _09658_/B _09658_/Y VGND VGND VPWR VPWR _10780_/X sky130_fd_sc_hd__o21a_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09439_ _09431_/A _09431_/B _09431_/X _09438_/X VGND VGND VPWR VPWR _09439_/X sky130_fd_sc_hd__a22o_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _13972_/A _12449_/B _12449_/Y VGND VGND VPWR VPWR _12450_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11401_ _11401_/A VGND VGND VPWR VPWR _11401_/Y sky130_fd_sc_hd__inv_2
X_14120_ _14120_/A VGND VGND VPWR VPWR _14120_/Y sky130_fd_sc_hd__inv_2
X_12381_ _12382_/A _12382_/B VGND VGND VPWR VPWR _12381_/X sky130_fd_sc_hd__and2_1
XFILLER_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11332_ _11331_/A _11331_/B _11331_/Y _10984_/X VGND VGND VPWR VPWR _12376_/A sky130_fd_sc_hd__o211a_1
XFILLER_125_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14051_ _15464_/A _14035_/B _14035_/X _14050_/X VGND VGND VPWR VPWR _14051_/X sky130_fd_sc_hd__o22a_1
X_11263_ _15443_/A _11179_/B _11179_/Y _11262_/X VGND VGND VPWR VPWR _11263_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11194_ _14057_/A VGND VGND VPWR VPWR _15449_/A sky130_fd_sc_hd__buf_1
XFILLER_79_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13002_ _12924_/A _13001_/Y _12924_/A _13001_/Y VGND VGND VPWR VPWR _13012_/B sky130_fd_sc_hd__a2bb2o_1
X_10214_ _10201_/Y _10212_/X _10213_/Y VGND VGND VPWR VPWR _10309_/B sky130_fd_sc_hd__o21ai_2
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10145_ _10147_/A VGND VGND VPWR VPWR _10240_/B sky130_fd_sc_hd__buf_1
XFILLER_121_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14953_ _14953_/A _14953_/B VGND VGND VPWR VPWR _14953_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10076_ _10075_/A _10075_/B _09700_/A _10075_/X VGND VGND VPWR VPWR _10076_/X sky130_fd_sc_hd__a22o_1
X_14884_ _14794_/A _14794_/B _14794_/A _14794_/B VGND VGND VPWR VPWR _14884_/X sky130_fd_sc_hd__a2bb2o_1
X_13904_ _15412_/A _13953_/B VGND VGND VPWR VPWR _13904_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13835_ _13754_/A _13834_/Y _13754_/A _13834_/Y VGND VGND VPWR VPWR _13837_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13766_ _13766_/A _13766_/B VGND VGND VPWR VPWR _13766_/X sky130_fd_sc_hd__or2_1
X_10978_ _12176_/A _11140_/B VGND VGND VPWR VPWR _10978_/Y sky130_fd_sc_hd__nand2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15505_ _15480_/X _15504_/X _15480_/X _15504_/X VGND VGND VPWR VPWR _15542_/B sky130_fd_sc_hd__a2bb2o_1
X_13697_ _13732_/A _13695_/X _13696_/X VGND VGND VPWR VPWR _13697_/X sky130_fd_sc_hd__o21a_1
X_12717_ _12691_/A _12691_/B _12691_/Y _12716_/X VGND VGND VPWR VPWR _12717_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12648_ _12495_/Y _12647_/X _12495_/Y _12647_/X VGND VGND VPWR VPWR _12649_/B sky130_fd_sc_hd__a2bb2oi_1
X_15436_ _15419_/X _15435_/Y _15419_/X _15435_/Y VGND VGND VPWR VPWR _15437_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12579_ _12579_/A VGND VGND VPWR VPWR _12579_/Y sky130_fd_sc_hd__inv_2
X_15367_ _15346_/X _15366_/X _15346_/X _15366_/X VGND VGND VPWR VPWR _15414_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14318_ _13437_/A _13437_/B _13437_/Y VGND VGND VPWR VPWR _14318_/X sky130_fd_sc_hd__o21a_1
X_15298_ _15281_/X _15297_/Y _15281_/X _15297_/Y VGND VGND VPWR VPWR _15349_/B sky130_fd_sc_hd__a2bb2o_1
X_14249_ _14371_/A _15885_/A VGND VGND VPWR VPWR _14249_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08810_ _10015_/A _08810_/B VGND VGND VPWR VPWR _08810_/Y sky130_fd_sc_hd__nor2_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09169_/A _09790_/A2 _09750_/Y _09789_/X VGND VGND VPWR VPWR _09793_/A sky130_fd_sc_hd__o22a_1
XFILLER_112_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08741_ _08710_/Y _08739_/Y _08740_/X VGND VGND VPWR VPWR _08742_/A sky130_fd_sc_hd__o21ai_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08672_ _09680_/A VGND VGND VPWR VPWR _10098_/A sky130_fd_sc_hd__inv_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09224_ _09224_/A VGND VGND VPWR VPWR _09224_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09155_ _09527_/B _09155_/B VGND VGND VPWR VPWR _09156_/B sky130_fd_sc_hd__or2_1
XFILLER_107_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09086_ _09769_/A VGND VGND VPWR VPWR _09424_/A sky130_fd_sc_hd__buf_1
XFILLER_107_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09988_ _09968_/Y _09986_/Y _09987_/Y VGND VGND VPWR VPWR _09990_/B sky130_fd_sc_hd__o21ai_2
X_08939_ _08942_/A _08942_/B VGND VGND VPWR VPWR _08939_/Y sky130_fd_sc_hd__nor2_1
X_11950_ _11903_/A _11949_/Y _11903_/A _11949_/Y VGND VGND VPWR VPWR _11972_/B sky130_fd_sc_hd__a2bb2o_1
X_10901_ _13184_/A _10912_/B VGND VGND VPWR VPWR _10901_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11881_ _11841_/X _11880_/Y _11841_/X _11880_/Y VGND VGND VPWR VPWR _11901_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13620_ _13620_/A VGND VGND VPWR VPWR _15137_/A sky130_fd_sc_hd__buf_1
X_10832_ _10964_/A _12082_/A VGND VGND VPWR VPWR _10832_/Y sky130_fd_sc_hd__nor2_1
X_10763_ _10763_/A _12606_/A VGND VGND VPWR VPWR _13753_/A sky130_fd_sc_hd__or2_1
X_13551_ _13551_/A _13551_/B VGND VGND VPWR VPWR _13552_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16270_ _16270_/A _16270_/B VGND VGND VPWR VPWR _16270_/Y sky130_fd_sc_hd__nand2_1
X_12502_ _12502_/A VGND VGND VPWR VPWR _12503_/A sky130_fd_sc_hd__buf_6
X_15221_ _15202_/A _15202_/B _15202_/Y _15220_/X VGND VGND VPWR VPWR _15221_/X sky130_fd_sc_hd__a2bb2o_1
X_13482_ _10296_/A _12702_/A _10325_/Y _13481_/X VGND VGND VPWR VPWR _13482_/X sky130_fd_sc_hd__o22a_1
X_10694_ _11992_/A VGND VGND VPWR VPWR _12693_/A sky130_fd_sc_hd__buf_1
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12433_ _12422_/A _12422_/B _12427_/X _12422_/Y _12432_/Y VGND VGND VPWR VPWR _12433_/X
+ sky130_fd_sc_hd__a32o_1
X_12364_ _12364_/A _12364_/B VGND VGND VPWR VPWR _12364_/Y sky130_fd_sc_hd__nor2_1
X_15152_ _15131_/A _15131_/B _15131_/Y _15151_/X VGND VGND VPWR VPWR _15152_/X sky130_fd_sc_hd__a2bb2o_1
X_14103_ _15458_/A _14027_/B _14027_/A _14027_/B VGND VGND VPWR VPWR _14103_/X sky130_fd_sc_hd__a2bb2o_1
X_15083_ _15027_/X _15082_/X _15027_/X _15082_/X VGND VGND VPWR VPWR _15084_/B sky130_fd_sc_hd__a2bb2o_1
X_11315_ _11311_/Y _12687_/A _11139_/X _11314_/Y VGND VGND VPWR VPWR _11315_/X sky130_fd_sc_hd__o22a_1
X_14034_ _13942_/X _14033_/Y _13942_/X _14033_/Y VGND VGND VPWR VPWR _14035_/B sky130_fd_sc_hd__a2bb2o_1
X_12295_ _13889_/A _12296_/B VGND VGND VPWR VPWR _12295_/X sky130_fd_sc_hd__and2_1
XFILLER_122_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11246_ _11246_/A VGND VGND VPWR VPWR _13935_/B sky130_fd_sc_hd__buf_1
XFILLER_122_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11177_ _11177_/A _11176_/X VGND VGND VPWR VPWR _11177_/X sky130_fd_sc_hd__or2b_1
X_15985_ _15984_/Y _15979_/X _15976_/Y VGND VGND VPWR VPWR _15985_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10128_ _10128_/A _10128_/B VGND VGND VPWR VPWR _10129_/B sky130_fd_sc_hd__or2_1
X_14936_ _12786_/A _12385_/B _12385_/Y _14839_/X VGND VGND VPWR VPWR _14936_/X sky130_fd_sc_hd__o2bb2a_1
X_10059_ _10059_/A _10059_/B VGND VGND VPWR VPWR _10059_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14867_ _15550_/A _14926_/B VGND VGND VPWR VPWR _14867_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14798_ _14798_/A _14798_/B VGND VGND VPWR VPWR _14798_/X sky130_fd_sc_hd__and2_1
XFILLER_90_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13818_ _13818_/A _13762_/X VGND VGND VPWR VPWR _13818_/X sky130_fd_sc_hd__or2b_1
XFILLER_23_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13749_ _13756_/A _13756_/B VGND VGND VPWR VPWR _13749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16468_ _08229_/A _16468_/D VGND VGND VPWR VPWR _16468_/Q sky130_fd_sc_hd__dfxtp_1
X_16399_ _16402_/B VGND VGND VPWR VPWR _16399_/Y sky130_fd_sc_hd__inv_2
X_15419_ _15362_/X _15417_/X _15438_/B VGND VGND VPWR VPWR _15419_/X sky130_fd_sc_hd__o21a_1
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09911_ _09908_/X _09911_/B VGND VGND VPWR VPWR _09913_/B sky130_fd_sc_hd__nand2b_1
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09842_ _09843_/A _09843_/B VGND VGND VPWR VPWR _10490_/A sky130_fd_sc_hd__and2_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A _09773_/B VGND VGND VPWR VPWR _09773_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08724_ _09228_/A _09458_/B VGND VGND VPWR VPWR _08724_/X sky130_fd_sc_hd__or2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08655_ _09799_/A VGND VGND VPWR VPWR _09684_/A sky130_fd_sc_hd__inv_2
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08586_ _08586_/A VGND VGND VPWR VPWR _08586_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09207_ _14011_/A VGND VGND VPWR VPWR _14061_/A sky130_fd_sc_hd__buf_1
XFILLER_22_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09138_ _09436_/A _09141_/B VGND VGND VPWR VPWR _09138_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11100_ _12261_/A VGND VGND VPWR VPWR _13712_/A sky130_fd_sc_hd__buf_1
X_09069_ _09069_/A _09069_/B VGND VGND VPWR VPWR _09070_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12080_ _12080_/A VGND VGND VPWR VPWR _12169_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_104_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11031_ _12847_/A VGND VGND VPWR VPWR _15072_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15770_ _15781_/B _15770_/B VGND VGND VPWR VPWR _16086_/A sky130_fd_sc_hd__or2_1
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12982_ _12935_/X _12981_/Y _12935_/X _12981_/Y VGND VGND VPWR VPWR _13023_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14721_ _14721_/A _14721_/B VGND VGND VPWR VPWR _14721_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11933_ _11987_/B _11932_/Y _11987_/B _11932_/Y VGND VGND VPWR VPWR _11985_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_45_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14652_ _14629_/Y _14650_/X _14651_/Y VGND VGND VPWR VPWR _14652_/X sky130_fd_sc_hd__o21a_1
X_11864_ _11921_/B _11863_/Y _11921_/B _11863_/Y VGND VGND VPWR VPWR _11917_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13603_ _13567_/A _13567_/B _13568_/A VGND VGND VPWR VPWR _13603_/Y sky130_fd_sc_hd__o21ai_1
X_10815_ _10814_/Y _10678_/X _10687_/Y VGND VGND VPWR VPWR _10815_/X sky130_fd_sc_hd__o21a_1
X_16322_ _16322_/A _16322_/B VGND VGND VPWR VPWR _16322_/Y sky130_fd_sc_hd__nand2_1
X_14583_ _14583_/A _14583_/B VGND VGND VPWR VPWR _14583_/Y sky130_fd_sc_hd__nand2_1
X_11795_ _11795_/A _11795_/B VGND VGND VPWR VPWR _11795_/X sky130_fd_sc_hd__or2_1
X_10746_ _11968_/A VGND VGND VPWR VPWR _13088_/A sky130_fd_sc_hd__buf_1
X_13534_ _15034_/A _13521_/B _13521_/Y _13533_/X VGND VGND VPWR VPWR _13534_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16253_ _16253_/A _16253_/B VGND VGND VPWR VPWR _16253_/Y sky130_fd_sc_hd__nand2_1
X_13465_ _13460_/Y _13464_/Y _13460_/Y _13464_/Y VGND VGND VPWR VPWR _13465_/X sky130_fd_sc_hd__a2bb2o_1
X_10677_ _11923_/A _10677_/B VGND VGND VPWR VPWR _10677_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16184_ _16192_/A _16184_/B VGND VGND VPWR VPWR _16262_/B sky130_fd_sc_hd__or2_1
X_15204_ _15149_/X _15203_/Y _15149_/X _15203_/Y VGND VGND VPWR VPWR _15205_/B sky130_fd_sc_hd__a2bb2o_1
X_12416_ _11614_/X _12425_/A _11614_/X _12425_/A VGND VGND VPWR VPWR _12429_/B sky130_fd_sc_hd__o2bb2a_1
X_13396_ _14097_/A VGND VGND VPWR VPWR _14100_/A sky130_fd_sc_hd__buf_1
X_15135_ _15078_/A _15078_/B _15078_/Y VGND VGND VPWR VPWR _15135_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12347_ _12343_/Y _12561_/A _12346_/Y VGND VGND VPWR VPWR _12351_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15066_ _15066_/A _15066_/B VGND VGND VPWR VPWR _15066_/Y sky130_fd_sc_hd__nand2_1
X_12278_ _12784_/A _12372_/A VGND VGND VPWR VPWR _12278_/Y sky130_fd_sc_hd__nor2_1
X_14017_ _14017_/A _14057_/B VGND VGND VPWR VPWR _14116_/A sky130_fd_sc_hd__and2_1
X_11229_ _11229_/A _11082_/X VGND VGND VPWR VPWR _11229_/X sky130_fd_sc_hd__or2b_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15968_ _15905_/X _15967_/Y _15905_/X _15967_/Y VGND VGND VPWR VPWR _15968_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15899_ _15865_/Y _15897_/X _15898_/Y VGND VGND VPWR VPWR _15899_/X sky130_fd_sc_hd__o21a_1
X_14919_ _14883_/Y _14917_/X _14918_/Y VGND VGND VPWR VPWR _14919_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08440_ _08440_/A VGND VGND VPWR VPWR _08440_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08371_ input15/X _08260_/B _08337_/B _08424_/A VGND VGND VPWR VPWR _08429_/A sky130_fd_sc_hd__o22a_1
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09825_ _09818_/A _09818_/B _09819_/B VGND VGND VPWR VPWR _09838_/A sky130_fd_sc_hd__a21bo_1
XFILLER_101_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09756_ _10085_/A VGND VGND VPWR VPWR _09995_/B sky130_fd_sc_hd__buf_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08707_ _09448_/B VGND VGND VPWR VPWR _08755_/A sky130_fd_sc_hd__inv_2
X_09687_ _09687_/A _09687_/B VGND VGND VPWR VPWR _09690_/B sky130_fd_sc_hd__or2_1
XFILLER_27_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08638_ _08483_/X _08388_/A _08483_/X _08388_/A VGND VGND VPWR VPWR _08639_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _09453_/B VGND VGND VPWR VPWR _08713_/B sky130_fd_sc_hd__inv_2
XFILLER_30_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10600_ _13620_/A _10529_/B _10529_/Y VGND VGND VPWR VPWR _10600_/Y sky130_fd_sc_hd__o21ai_1
X_11580_ _11579_/A _11579_/B _11579_/Y _09392_/X VGND VGND VPWR VPWR _13133_/A sky130_fd_sc_hd__o211a_1
XFILLER_10_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10531_ _11844_/A _10531_/B VGND VGND VPWR VPWR _10531_/Y sky130_fd_sc_hd__nand2_1
X_13250_ _14730_/A _13285_/B VGND VGND VPWR VPWR _13250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12201_ _13893_/A _12202_/B VGND VGND VPWR VPWR _12201_/X sky130_fd_sc_hd__and2_1
X_10462_ _10462_/A VGND VGND VPWR VPWR _10976_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13181_ _13096_/X _13180_/Y _13096_/A _13180_/Y VGND VGND VPWR VPWR _13182_/B sky130_fd_sc_hd__a2bb2o_1
X_10393_ _10245_/A _09306_/B _09306_/Y VGND VGND VPWR VPWR _10394_/A sky130_fd_sc_hd__o21ai_1
X_12132_ _12050_/X _12131_/Y _12050_/X _12131_/Y VGND VGND VPWR VPWR _12139_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12063_ _12063_/A _12063_/B VGND VGND VPWR VPWR _12063_/Y sky130_fd_sc_hd__nand2_1
X_11014_ _10923_/X _11013_/X _10923_/X _11013_/X VGND VGND VPWR VPWR _11092_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15822_ _15712_/X _15820_/X _16142_/B VGND VGND VPWR VPWR _15822_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15753_ _15675_/A _15675_/B _15675_/Y VGND VGND VPWR VPWR _15753_/Y sky130_fd_sc_hd__o21ai_1
X_12965_ _14676_/A _12944_/B _12944_/Y VGND VGND VPWR VPWR _12965_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14704_ _14730_/A _14730_/B VGND VGND VPWR VPWR _14796_/A sky130_fd_sc_hd__and2_1
XFILLER_73_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11916_ _11916_/A _11916_/B VGND VGND VPWR VPWR _11916_/X sky130_fd_sc_hd__or2_1
XFILLER_45_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15684_ _15592_/Y _15682_/X _15683_/Y VGND VGND VPWR VPWR _15684_/X sky130_fd_sc_hd__o21a_1
X_12896_ _14466_/A _12934_/B VGND VGND VPWR VPWR _12896_/Y sky130_fd_sc_hd__nor2_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14575_/A _14575_/B _14575_/Y VGND VGND VPWR VPWR _14635_/Y sky130_fd_sc_hd__o21ai_1
X_11847_ _11821_/Y _11845_/X _11846_/Y VGND VGND VPWR VPWR _11847_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _15272_/A _14573_/B VGND VGND VPWR VPWR _14566_/Y sky130_fd_sc_hd__nor2_1
X_11778_ _11778_/A _11778_/B VGND VGND VPWR VPWR _11778_/X sky130_fd_sc_hd__and2_1
XFILLER_13_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16305_ _16322_/A _16322_/B VGND VGND VPWR VPWR _16305_/Y sky130_fd_sc_hd__nor2_1
X_10729_ _11972_/A VGND VGND VPWR VPWR _13078_/A sky130_fd_sc_hd__buf_1
X_13517_ _10475_/X _13484_/X _10475_/X _13484_/X VGND VGND VPWR VPWR _13518_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16236_ _16089_/A _15790_/B _15790_/Y VGND VGND VPWR VPWR _16236_/X sky130_fd_sc_hd__o21a_1
X_14497_ _14460_/A _14460_/B _14460_/Y VGND VGND VPWR VPWR _14497_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13448_ _13377_/Y _13446_/X _13447_/Y VGND VGND VPWR VPWR _13448_/X sky130_fd_sc_hd__o21a_1
X_16167_ _15814_/X _16166_/X _15814_/X _16166_/X VGND VGND VPWR VPWR _16168_/B sky130_fd_sc_hd__a2bb2o_1
X_13379_ _13369_/X _13378_/X _13369_/X _13378_/X VGND VGND VPWR VPWR _13445_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16098_ _16033_/X _16097_/Y _16033_/X _16097_/Y VGND VGND VPWR VPWR _16098_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15118_ _15096_/X _15117_/Y _15096_/X _15117_/Y VGND VGND VPWR VPWR _15119_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15049_ _12276_/Y _15048_/X _12276_/Y _15048_/X VGND VGND VPWR VPWR _15051_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09610_ _09496_/A _09496_/B _09496_/Y VGND VGND VPWR VPWR _09610_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09541_ _09541_/A _09541_/B VGND VGND VPWR VPWR _09629_/B sky130_fd_sc_hd__or2_1
XFILLER_64_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09472_ _10011_/A _09472_/B VGND VGND VPWR VPWR _09472_/X sky130_fd_sc_hd__or2_1
X_08423_ _09217_/B _08417_/Y _09249_/A VGND VGND VPWR VPWR _08423_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08354_ _08354_/A VGND VGND VPWR VPWR _08354_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08285_ input27/X _08363_/B _08364_/A _08384_/A VGND VGND VPWR VPWR _08355_/A sky130_fd_sc_hd__o22a_1
XFILLER_20_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09808_ _09808_/A VGND VGND VPWR VPWR _09826_/A sky130_fd_sc_hd__inv_2
XFILLER_74_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09739_ _09739_/A _09739_/B VGND VGND VPWR VPWR _09742_/A sky130_fd_sc_hd__or2_1
XFILLER_55_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12750_ _12712_/X _12749_/X _12712_/X _12749_/X VGND VGND VPWR VPWR _12770_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _12454_/A VGND VGND VPWR VPWR _13978_/A sky130_fd_sc_hd__clkbuf_2
X_12681_ _12428_/A _12680_/B _12680_/Y VGND VGND VPWR VPWR _12681_/X sky130_fd_sc_hd__a21o_1
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/A _14420_/B VGND VGND VPWR VPWR _14420_/Y sky130_fd_sc_hd__nor2_1
X_11632_ _11632_/A _11632_/B VGND VGND VPWR VPWR _11632_/Y sky130_fd_sc_hd__nor2_1
X_14351_ _13414_/Y _14350_/X _13414_/Y _14350_/X VGND VGND VPWR VPWR _14352_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_128_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13302_ _13302_/A VGND VGND VPWR VPWR _13302_/Y sky130_fd_sc_hd__inv_2
X_11563_ _11474_/X _11562_/X _11474_/X _11562_/X VGND VGND VPWR VPWR _11564_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14282_ _14285_/A _15908_/A VGND VGND VPWR VPWR _14282_/X sky130_fd_sc_hd__and2_1
X_11494_ _11494_/A VGND VGND VPWR VPWR _11494_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10514_ _09829_/A _09829_/B _09830_/A VGND VGND VPWR VPWR _10514_/Y sky130_fd_sc_hd__o21ai_1
X_16021_ _15949_/X _16020_/Y _15949_/X _16020_/Y VGND VGND VPWR VPWR _16032_/B sky130_fd_sc_hd__a2bb2o_1
X_13233_ _13198_/A _13198_/B _13198_/Y VGND VGND VPWR VPWR _13233_/Y sky130_fd_sc_hd__o21ai_1
X_10445_ _10445_/A VGND VGND VPWR VPWR _10959_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13164_ _13110_/X _13163_/Y _13110_/X _13163_/Y VGND VGND VPWR VPWR _13192_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12115_ _13905_/A _12151_/B VGND VGND VPWR VPWR _12212_/A sky130_fd_sc_hd__and2_1
X_10376_ _10376_/A VGND VGND VPWR VPWR _10376_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13095_ _14563_/A _13103_/B VGND VGND VPWR VPWR _13095_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12046_ _10768_/A _11964_/B _10768_/A _11964_/B VGND VGND VPWR VPWR _12046_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15805_ _16104_/A _15805_/B VGND VGND VPWR VPWR _15805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13997_ _13997_/A VGND VGND VPWR VPWR _13997_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15736_ _15680_/X _15735_/Y _15680_/X _15735_/Y VGND VGND VPWR VPWR _15813_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12948_ _12948_/A VGND VGND VPWR VPWR _14944_/A sky130_fd_sc_hd__buf_1
X_15667_ _15667_/A _15667_/B VGND VGND VPWR VPWR _15788_/B sky130_fd_sc_hd__or2_1
XFILLER_61_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12879_ _12854_/X _12878_/Y _12854_/X _12878_/Y VGND VGND VPWR VPWR _12942_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14618_ _14618_/A VGND VGND VPWR VPWR _15341_/A sky130_fd_sc_hd__buf_1
XFILLER_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15598_ _14390_/X _15597_/Y _14390_/X _15597_/Y VGND VGND VPWR VPWR _15681_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14549_ _14516_/X _14548_/X _14516_/X _14548_/X VGND VGND VPWR VPWR _14581_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16219_ _16217_/A _16218_/A _16217_/Y _16218_/Y _15832_/A VGND VGND VPWR VPWR _16253_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08972_ _08972_/A _08972_/B VGND VGND VPWR VPWR _11387_/B sky130_fd_sc_hd__or2_1
XFILLER_96_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09524_ _09561_/A _09561_/B VGND VGND VPWR VPWR _09567_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09455_ _09494_/A _09455_/B VGND VGND VPWR VPWR _09455_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08406_ _08944_/A VGND VGND VPWR VPWR _09459_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09386_ _09430_/B _09370_/B _09370_/X _11476_/A VGND VGND VPWR VPWR _11579_/A sky130_fd_sc_hd__a22o_1
X_08337_ _08337_/A _08337_/B VGND VGND VPWR VPWR _08338_/A sky130_fd_sc_hd__or2_1
X_08268_ input28/X VGND VGND VPWR VPWR _08269_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_20_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10230_ _10230_/A _10230_/B VGND VGND VPWR VPWR _10231_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10161_ _10163_/A VGND VGND VPWR VPWR _10244_/B sky130_fd_sc_hd__buf_1
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10092_ _10007_/X _10091_/X _10007_/X _10091_/X VGND VGND VPWR VPWR _10215_/A sky130_fd_sc_hd__a2bb2o_4
X_13920_ _15404_/A _13945_/B VGND VGND VPWR VPWR _13920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13851_ _14614_/A _13851_/B VGND VGND VPWR VPWR _13851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10994_ _12097_/A _11122_/B VGND VGND VPWR VPWR _10994_/Y sky130_fd_sc_hd__nand2_1
X_12802_ _12855_/A _12855_/B VGND VGND VPWR VPWR _12802_/Y sky130_fd_sc_hd__nor2_1
X_13782_ _12857_/A _13712_/B _13781_/Y _13709_/X VGND VGND VPWR VPWR _13782_/X sky130_fd_sc_hd__o22a_1
XFILLER_43_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15521_ _15524_/A _15524_/B VGND VGND VPWR VPWR _15521_/Y sky130_fd_sc_hd__nor2_1
X_12733_ _12782_/A _12782_/B VGND VGND VPWR VPWR _12733_/Y sky130_fd_sc_hd__nor2_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _15452_/A _15452_/B VGND VGND VPWR VPWR _15452_/X sky130_fd_sc_hd__and2_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14403_ _14296_/Y _14401_/X _14402_/Y VGND VGND VPWR VPWR _14403_/X sky130_fd_sc_hd__o21a_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _10556_/Y _12663_/Y _10464_/Y VGND VGND VPWR VPWR _12665_/A sky130_fd_sc_hd__o21ai_1
XFILLER_129_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12595_ _12595_/A VGND VGND VPWR VPWR _12595_/Y sky130_fd_sc_hd__inv_2
X_15383_ _15404_/A _15404_/B VGND VGND VPWR VPWR _15459_/A sky130_fd_sc_hd__and2_1
X_11615_ _11615_/A _11615_/B VGND VGND VPWR VPWR _11615_/Y sky130_fd_sc_hd__nor2_1
X_14334_ _14334_/A _14334_/B VGND VGND VPWR VPWR _15956_/A sky130_fd_sc_hd__or2_1
X_11546_ _12390_/A _11641_/B VGND VGND VPWR VPWR _11546_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14265_ _15866_/A _14265_/B VGND VGND VPWR VPWR _14265_/Y sky130_fd_sc_hd__nand2_1
X_16004_ _16044_/A _16044_/B VGND VGND VPWR VPWR _16004_/Y sky130_fd_sc_hd__nor2_1
X_13216_ _15054_/A VGND VGND VPWR VPWR _14754_/A sky130_fd_sc_hd__inv_2
X_11477_ _11476_/A _11476_/B _11476_/Y _09392_/X VGND VGND VPWR VPWR _12442_/A sky130_fd_sc_hd__o211a_1
XFILLER_7_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14196_ _12629_/X _14195_/X _12629_/X _14195_/X VGND VGND VPWR VPWR _14268_/B sky130_fd_sc_hd__a2bb2o_1
X_10428_ _10625_/A VGND VGND VPWR VPWR _10428_/X sky130_fd_sc_hd__buf_1
XFILLER_124_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13147_ _13204_/A _13204_/B VGND VGND VPWR VPWR _13147_/Y sky130_fd_sc_hd__nor2_1
X_10359_ _13527_/A _10328_/B _10328_/X _10358_/X VGND VGND VPWR VPWR _10359_/X sky130_fd_sc_hd__o22a_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13078_ _13078_/A VGND VGND VPWR VPWR _13762_/A sky130_fd_sc_hd__inv_2
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _12057_/A VGND VGND VPWR VPWR _13190_/A sky130_fd_sc_hd__buf_1
XFILLER_78_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15719_ _15548_/A _14924_/B _14924_/Y VGND VGND VPWR VPWR _15719_/X sky130_fd_sc_hd__o21a_1
X_09240_ _08623_/A _09802_/A _09224_/Y _09239_/Y VGND VGND VPWR VPWR _09240_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09171_ _10009_/B _09166_/B _09167_/B VGND VGND VPWR VPWR _09754_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08955_ _08955_/A VGND VGND VPWR VPWR _08955_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08886_ _08886_/A _08886_/B VGND VGND VPWR VPWR _08886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09507_ _09502_/A _09502_/B _09502_/Y _09506_/X VGND VGND VPWR VPWR _09507_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09438_ _09432_/A _09432_/B _09432_/X _11107_/A VGND VGND VPWR VPWR _09438_/X sky130_fd_sc_hd__a22o_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09369_ _10238_/A VGND VGND VPWR VPWR _09370_/B sky130_fd_sc_hd__buf_1
X_12380_ _11533_/Y _12379_/X _11533_/Y _12379_/X VGND VGND VPWR VPWR _12382_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11400_ _08960_/A _08960_/B _08960_/Y VGND VGND VPWR VPWR _11401_/A sky130_fd_sc_hd__o21ai_1
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11331_ _11331_/A _11331_/B VGND VGND VPWR VPWR _11331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14050_ _13344_/A _14038_/B _14038_/X _14049_/X VGND VGND VPWR VPWR _14050_/X sky130_fd_sc_hd__o22a_1
X_11262_ _15446_/A _11188_/B _11188_/Y _11261_/X VGND VGND VPWR VPWR _11262_/X sky130_fd_sc_hd__a2bb2o_1
X_11193_ _14017_/A VGND VGND VPWR VPWR _14057_/A sky130_fd_sc_hd__buf_1
XFILLER_97_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13001_ _14458_/A _12926_/B _12926_/Y VGND VGND VPWR VPWR _13001_/Y sky130_fd_sc_hd__o21ai_1
X_10213_ _10213_/A _10213_/B VGND VGND VPWR VPWR _10213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10144_ _10118_/A _10118_/B _10119_/A VGND VGND VPWR VPWR _10147_/A sky130_fd_sc_hd__a21bo_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14952_ _14976_/A _14976_/B _14951_/Y VGND VGND VPWR VPWR _14952_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10075_ _10075_/A _10075_/B VGND VGND VPWR VPWR _10075_/X sky130_fd_sc_hd__or2_1
X_14883_ _15542_/A _14918_/B VGND VGND VPWR VPWR _14883_/Y sky130_fd_sc_hd__nor2_1
X_13903_ _13852_/X _13902_/Y _13852_/X _13902_/Y VGND VGND VPWR VPWR _13953_/B sky130_fd_sc_hd__a2bb2o_1
X_13834_ _13752_/A _13752_/B _13752_/Y VGND VGND VPWR VPWR _13834_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13765_ _13815_/A _13763_/X _13764_/X VGND VGND VPWR VPWR _13765_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10977_ _10975_/A _10974_/Y _10975_/Y _10974_/A _11529_/A VGND VGND VPWR VPWR _11140_/B
+ sky130_fd_sc_hd__a221o_1
X_15504_ _15452_/A _15452_/B _15452_/A _15452_/B VGND VGND VPWR VPWR _15504_/X sky130_fd_sc_hd__a2bb2o_1
X_13696_ _13696_/A _13696_/B VGND VGND VPWR VPWR _13696_/X sky130_fd_sc_hd__or2_1
X_12716_ _12693_/A _12693_/B _12693_/Y _12715_/X VGND VGND VPWR VPWR _12716_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12647_ _14984_/A _12496_/B _12496_/Y VGND VGND VPWR VPWR _12647_/X sky130_fd_sc_hd__o21a_1
X_15435_ _15359_/X _15435_/B VGND VGND VPWR VPWR _15435_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_129_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15366_ _15366_/A _15347_/X VGND VGND VPWR VPWR _15366_/X sky130_fd_sc_hd__or2b_1
X_12578_ _14910_/A _11437_/B _11437_/Y VGND VGND VPWR VPWR _12579_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14317_ _15962_/A _14391_/B VGND VGND VPWR VPWR _14317_/X sky130_fd_sc_hd__and2_1
X_15297_ _14745_/A _15240_/B _15240_/Y VGND VGND VPWR VPWR _15297_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11529_ _11529_/A _11529_/B VGND VGND VPWR VPWR _11615_/B sky130_fd_sc_hd__or2_1
X_14248_ _14371_/B _14248_/B VGND VGND VPWR VPWR _15885_/A sky130_fd_sc_hd__nor2_1
X_14179_ _15906_/A _14277_/B VGND VGND VPWR VPWR _14179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08740_ _10010_/A _09527_/A VGND VGND VPWR VPWR _08740_/X sky130_fd_sc_hd__or2_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08671_ _08671_/A _08929_/A VGND VGND VPWR VPWR _09680_/A sky130_fd_sc_hd__or2_1
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09223_ _09547_/A _09693_/A VGND VGND VPWR VPWR _09224_/A sky130_fd_sc_hd__or2_1
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09154_ _09154_/A VGND VGND VPWR VPWR _09527_/B sky130_fd_sc_hd__inv_2
X_09085_ _10014_/B _09075_/B _09076_/B VGND VGND VPWR VPWR _09769_/A sky130_fd_sc_hd__a21bo_1
XFILLER_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09987_ _09987_/A _09987_/B VGND VGND VPWR VPWR _09987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08938_ _08936_/Y _08937_/X _08936_/Y _08937_/X VGND VGND VPWR VPWR _08942_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08869_ _08753_/Y _08868_/Y _08753_/Y _08868_/Y VGND VGND VPWR VPWR _08986_/B sky130_fd_sc_hd__o2bb2a_1
X_10900_ _10770_/X _10899_/X _10770_/X _10899_/X VGND VGND VPWR VPWR _10912_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11880_ _11842_/A _11842_/B _11842_/Y VGND VGND VPWR VPWR _11880_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10831_ _12082_/A VGND VGND VPWR VPWR _12691_/A sky130_fd_sc_hd__buf_1
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10762_ _10768_/A _10769_/B VGND VGND VPWR VPWR _10904_/A sky130_fd_sc_hd__and2_1
X_13550_ _13535_/X _13549_/Y _13535_/X _13549_/Y VGND VGND VPWR VPWR _13551_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12501_ _12501_/A VGND VGND VPWR VPWR _12502_/A sky130_fd_sc_hd__buf_6
X_13481_ _11734_/A _10294_/Y _10335_/Y _13480_/Y VGND VGND VPWR VPWR _13481_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15220_ _15205_/A _15205_/B _15205_/Y _15219_/X VGND VGND VPWR VPWR _15220_/X sky130_fd_sc_hd__a2bb2o_1
X_12432_ _12432_/A VGND VGND VPWR VPWR _12432_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10693_ _10692_/A _10692_/B _10692_/Y _10984_/A VGND VGND VPWR VPWR _11992_/A sky130_fd_sc_hd__o211a_1
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12363_ _12362_/Y _12255_/X _12289_/Y VGND VGND VPWR VPWR _12363_/Y sky130_fd_sc_hd__o21ai_1
X_15151_ _15134_/A _15134_/B _15134_/Y _15150_/X VGND VGND VPWR VPWR _15151_/X sky130_fd_sc_hd__a2bb2o_1
X_14102_ _14102_/A _14105_/B VGND VGND VPWR VPWR _14102_/Y sky130_fd_sc_hd__nor2_1
X_12294_ _12252_/X _12293_/Y _12252_/X _12293_/Y VGND VGND VPWR VPWR _12296_/B sky130_fd_sc_hd__a2bb2o_1
X_15082_ _15082_/A _15028_/X VGND VGND VPWR VPWR _15082_/X sky130_fd_sc_hd__or2b_1
X_11314_ _11314_/A _12181_/A VGND VGND VPWR VPWR _11314_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11245_ _11245_/A _11413_/B VGND VGND VPWR VPWR _14047_/A sky130_fd_sc_hd__or2_1
X_14033_ _15402_/A _13943_/B _13943_/Y VGND VGND VPWR VPWR _14033_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11176_ _13893_/A _11176_/B VGND VGND VPWR VPWR _11176_/X sky130_fd_sc_hd__or2_1
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15984_ _15984_/A _15984_/B VGND VGND VPWR VPWR _15984_/Y sky130_fd_sc_hd__nor2_1
X_10127_ _10127_/A _10127_/B VGND VGND VPWR VPWR _10128_/B sky130_fd_sc_hd__or2_1
X_14935_ _14835_/X _14849_/A _14848_/X VGND VGND VPWR VPWR _14935_/X sky130_fd_sc_hd__o21a_1
X_10058_ _10019_/X _10057_/Y _10019_/X _10057_/Y VGND VGND VPWR VPWR _10059_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14866_ _14826_/X _14865_/X _14826_/X _14865_/X VGND VGND VPWR VPWR _14926_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14797_ _14729_/X _14796_/X _14729_/X _14796_/X VGND VGND VPWR VPWR _14798_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13817_ _14622_/A _13847_/B VGND VGND VPWR VPWR _13817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13748_ _13685_/A _13747_/Y _13685_/A _13747_/Y VGND VGND VPWR VPWR _13756_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16467_ _08229_/A _16467_/D VGND VGND VPWR VPWR _16467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13679_ _14500_/A _13686_/B VGND VGND VPWR VPWR _13679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16398_ _16407_/B VGND VGND VPWR VPWR _16398_/Y sky130_fd_sc_hd__inv_2
X_15418_ _15418_/A _15418_/B VGND VGND VPWR VPWR _15438_/B sky130_fd_sc_hd__or2_1
XFILLER_117_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15349_ _15349_/A _15349_/B VGND VGND VPWR VPWR _15349_/X sky130_fd_sc_hd__or2_1
XFILLER_8_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09910_ _09908_/A _09908_/B _09909_/Y VGND VGND VPWR VPWR _09911_/B sky130_fd_sc_hd__o21ai_1
XFILLER_125_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09841_ _09838_/A _09838_/B _09839_/Y _10499_/A VGND VGND VPWR VPWR _09843_/B sky130_fd_sc_hd__o22a_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09773_/A _09773_/B VGND VGND VPWR VPWR _09772_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08723_ _08843_/A _09459_/B _08719_/Y _08722_/X VGND VGND VPWR VPWR _08723_/X sky130_fd_sc_hd__o22a_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ _08843_/A _09006_/A VGND VGND VPWR VPWR _09799_/A sky130_fd_sc_hd__or2_1
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08585_ _09467_/B _10115_/B VGND VGND VPWR VPWR _08586_/A sky130_fd_sc_hd__or2_1
XFILLER_81_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09206_ _13368_/A VGND VGND VPWR VPWR _14011_/A sky130_fd_sc_hd__inv_2
XFILLER_50_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09137_ _09133_/Y _09135_/Y _09136_/Y VGND VGND VPWR VPWR _09141_/B sky130_fd_sc_hd__o21ai_1
X_09068_ _10102_/A _09627_/A VGND VGND VPWR VPWR _09069_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11030_ _13555_/A VGND VGND VPWR VPWR _12847_/A sky130_fd_sc_hd__buf_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12981_ _14468_/A _12936_/B _12936_/Y VGND VGND VPWR VPWR _12981_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14720_ _14721_/A _14721_/B VGND VGND VPWR VPWR _14720_/Y sky130_fd_sc_hd__nor2_1
X_11932_ _12776_/A _11988_/A _11931_/Y VGND VGND VPWR VPWR _11932_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14651_ _15337_/A _14651_/B VGND VGND VPWR VPWR _14651_/Y sky130_fd_sc_hd__nand2_1
X_11863_ _11861_/X _11863_/B VGND VGND VPWR VPWR _11863_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13602_ _13605_/A VGND VGND VPWR VPWR _15140_/A sky130_fd_sc_hd__buf_1
XFILLER_60_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10814_ _11994_/A _10814_/B VGND VGND VPWR VPWR _10814_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16321_ _16308_/Y _16319_/X _16320_/Y VGND VGND VPWR VPWR _16321_/X sky130_fd_sc_hd__o21a_1
X_14582_ _14550_/Y _14580_/X _14581_/Y VGND VGND VPWR VPWR _14582_/X sky130_fd_sc_hd__o21a_1
X_11794_ _11794_/A _11794_/B VGND VGND VPWR VPWR _11794_/X sky130_fd_sc_hd__and2_1
XFILLER_13_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13533_ _15032_/A _13524_/B _13524_/Y _13532_/X VGND VGND VPWR VPWR _13533_/X sky130_fd_sc_hd__a2bb2o_1
X_10745_ _10743_/A _10744_/A _10743_/Y _10744_/Y _09672_/A VGND VGND VPWR VPWR _11968_/A
+ sky130_fd_sc_hd__a221o_2
X_16252_ _16231_/Y _16250_/X _16251_/Y VGND VGND VPWR VPWR _16252_/X sky130_fd_sc_hd__o21a_1
X_13464_ _13461_/Y _13463_/X _13461_/Y _13463_/X VGND VGND VPWR VPWR _13464_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10676_ _10673_/Y _12695_/A _10555_/X _10675_/Y VGND VGND VPWR VPWR _10676_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16183_ _15810_/X _16182_/X _15810_/X _16182_/X VGND VGND VPWR VPWR _16184_/B sky130_fd_sc_hd__a2bb2o_1
X_13395_ _13395_/A VGND VGND VPWR VPWR _14097_/A sky130_fd_sc_hd__inv_2
X_15203_ _15137_/A _15137_/B _15137_/Y VGND VGND VPWR VPWR _15203_/Y sky130_fd_sc_hd__o21ai_1
X_12415_ _11615_/A _11531_/B _12379_/X VGND VGND VPWR VPWR _12425_/A sky130_fd_sc_hd__o21ai_1
X_12346_ _12346_/A _12346_/B VGND VGND VPWR VPWR _12346_/Y sky130_fd_sc_hd__nand2_1
X_15134_ _15134_/A _15134_/B VGND VGND VPWR VPWR _15134_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15065_ _15039_/X _15064_/X _15039_/X _15064_/X VGND VGND VPWR VPWR _15066_/B sky130_fd_sc_hd__a2bb2o_1
X_12277_ _12376_/B _12276_/Y _12376_/B _12276_/Y VGND VGND VPWR VPWR _12372_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11228_ _14032_/A VGND VGND VPWR VPWR _14035_/A sky130_fd_sc_hd__buf_1
X_14016_ _13952_/X _14015_/Y _13952_/X _14015_/Y VGND VGND VPWR VPWR _14057_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11159_ _11139_/X _11158_/X _11139_/X _11158_/X VGND VGND VPWR VPWR _11306_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15967_ _15906_/A _15906_/B _15906_/Y VGND VGND VPWR VPWR _15967_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15898_ _15898_/A _15898_/B VGND VGND VPWR VPWR _15898_/Y sky130_fd_sc_hd__nand2_1
X_14918_ _15542_/A _14918_/B VGND VGND VPWR VPWR _14918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14849_ _14849_/A _14848_/X VGND VGND VPWR VPWR _14849_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08370_ _08263_/A input14/X _08342_/B _08418_/A VGND VGND VPWR VPWR _08424_/A sky130_fd_sc_hd__o22a_1
XFILLER_32_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09824_ _09819_/A _09819_/B _09820_/B VGND VGND VPWR VPWR _09843_/A sky130_fd_sc_hd__a21bo_1
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09742_/A _09742_/B _09745_/A VGND VGND VPWR VPWR _10085_/A sky130_fd_sc_hd__a21bo_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08706_ _09340_/A _08706_/B VGND VGND VPWR VPWR _08749_/A sky130_fd_sc_hd__or2_2
X_09686_ _09686_/A _09686_/B VGND VGND VPWR VPWR _09689_/A sky130_fd_sc_hd__or2_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _08637_/A VGND VGND VPWR VPWR _08637_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08568_ _08567_/X _08433_/X _08567_/X _08433_/X VGND VGND VPWR VPWR _08571_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08499_ _08650_/A VGND VGND VPWR VPWR _08589_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10530_ _10496_/Y _10528_/X _10529_/Y VGND VGND VPWR VPWR _10530_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10461_ _10461_/A VGND VGND VPWR VPWR _10461_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12200_ _12158_/X _12199_/Y _12158_/X _12199_/Y VGND VGND VPWR VPWR _12202_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13180_ _14567_/A _13101_/B _13101_/Y VGND VGND VPWR VPWR _13180_/Y sky130_fd_sc_hd__o21ai_1
X_10392_ _11773_/A _10392_/B VGND VGND VPWR VPWR _10392_/X sky130_fd_sc_hd__and2_1
XFILLER_123_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12131_ _13828_/A _12051_/B _12051_/Y VGND VGND VPWR VPWR _12131_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12062_ _12024_/Y _12060_/X _12061_/Y VGND VGND VPWR VPWR _12062_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11013_ _11013_/A _10925_/X VGND VGND VPWR VPWR _11013_/X sky130_fd_sc_hd__or2b_1
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15821_ _16123_/A _15821_/B VGND VGND VPWR VPWR _16142_/B sky130_fd_sc_hd__or2_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15752_ _15752_/A _15752_/B VGND VGND VPWR VPWR _16106_/A sky130_fd_sc_hd__nor2_1
X_12964_ _13719_/A VGND VGND VPWR VPWR _14668_/A sky130_fd_sc_hd__inv_2
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14703_ _14652_/X _14702_/Y _14652_/X _14702_/Y VGND VGND VPWR VPWR _14730_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11915_ _13551_/A _11914_/B _11914_/X _11849_/X VGND VGND VPWR VPWR _11915_/X sky130_fd_sc_hd__o22a_1
X_15683_ _15683_/A _15683_/B VGND VGND VPWR VPWR _15683_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12895_ _12846_/X _12894_/Y _12846_/X _12894_/Y VGND VGND VPWR VPWR _12934_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _14634_/A VGND VGND VPWR VPWR _15333_/A sky130_fd_sc_hd__buf_1
X_11846_ _11846_/A _11846_/B VGND VGND VPWR VPWR _11846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _14508_/X _14564_/X _14508_/X _14564_/X VGND VGND VPWR VPWR _14573_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11777_ _11744_/B _11776_/Y _11744_/B _11776_/Y VGND VGND VPWR VPWR _11778_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16304_ _16254_/X _16303_/Y _16254_/X _16303_/Y VGND VGND VPWR VPWR _16322_/B sky130_fd_sc_hd__o2bb2a_1
X_13516_ _13518_/A VGND VGND VPWR VPWR _15036_/A sky130_fd_sc_hd__buf_1
X_10728_ _10726_/A _10727_/A _10726_/Y _10727_/Y _09672_/A VGND VGND VPWR VPWR _11972_/A
+ sky130_fd_sc_hd__a221o_2
X_16235_ _16233_/A _16234_/A _16233_/Y _16234_/Y _16243_/A VGND VGND VPWR VPWR _16249_/A
+ sky130_fd_sc_hd__a221o_1
X_14496_ _14496_/A VGND VGND VPWR VPWR _15208_/A sky130_fd_sc_hd__buf_1
XFILLER_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13447_ _13447_/A _13447_/B VGND VGND VPWR VPWR _13447_/Y sky130_fd_sc_hd__nand2_1
X_10659_ _12938_/A VGND VGND VPWR VPWR _11936_/A sky130_fd_sc_hd__inv_2
X_16166_ _16114_/A _15815_/B _15815_/Y VGND VGND VPWR VPWR _16166_/X sky130_fd_sc_hd__o21a_1
X_13378_ _13378_/A _13370_/X VGND VGND VPWR VPWR _13378_/X sky130_fd_sc_hd__or2b_1
XFILLER_127_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16097_ _16034_/A _16034_/B _16034_/Y VGND VGND VPWR VPWR _16097_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12329_ _12229_/A _12229_/B _12229_/Y VGND VGND VPWR VPWR _12329_/Y sky130_fd_sc_hd__o21ai_1
X_15117_ _15060_/A _15060_/B _15060_/Y VGND VGND VPWR VPWR _15117_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15048_ _12182_/A _15006_/X _12181_/X VGND VGND VPWR VPWR _15048_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09540_ _09540_/A _09540_/B VGND VGND VPWR VPWR _09540_/X sky130_fd_sc_hd__or2_1
XFILLER_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09471_ _09452_/Y _09469_/X _09470_/X VGND VGND VPWR VPWR _09471_/X sky130_fd_sc_hd__o21a_1
X_08422_ _08715_/A VGND VGND VPWR VPWR _09249_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08353_ _08353_/A _08353_/B VGND VGND VPWR VPWR _08354_/A sky130_fd_sc_hd__or2_1
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08284_ input26/X _08357_/B _08387_/A _08389_/A VGND VGND VPWR VPWR _08384_/A sky130_fd_sc_hd__o22a_1
XFILLER_20_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09807_ _08852_/A _08721_/B _09817_/A VGND VGND VPWR VPWR _09808_/A sky130_fd_sc_hd__o21ai_1
X_09738_ _08546_/A _09740_/B _08546_/A _09740_/B VGND VGND VPWR VPWR _09739_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09669_ _09562_/Y _09668_/Y _09562_/Y _09668_/Y VGND VGND VPWR VPWR _09669_/X sky130_fd_sc_hd__a2bb2o_2
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11640_/A _11642_/X _11639_/X VGND VGND VPWR VPWR _11700_/X sky130_fd_sc_hd__o21a_1
X_12680_ _12680_/A _12680_/B VGND VGND VPWR VPWR _12680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11628_/Y _11630_/X _11628_/Y _11630_/X VGND VGND VPWR VPWR _11632_/B sky130_fd_sc_hd__o2bb2a_1
X_14350_ _13412_/X _14350_/B VGND VGND VPWR VPWR _14350_/X sky130_fd_sc_hd__and2b_1
X_11562_ _11562_/A _11561_/X VGND VGND VPWR VPWR _11562_/X sky130_fd_sc_hd__or2b_1
XFILLER_11_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13301_ _13225_/Y _13299_/Y _13300_/Y VGND VGND VPWR VPWR _13302_/A sky130_fd_sc_hd__o21ai_1
X_10513_ _15143_/A _10525_/B VGND VGND VPWR VPWR _10513_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14281_ _14281_/A _14281_/B VGND VGND VPWR VPWR _15908_/A sky130_fd_sc_hd__or2_1
X_11493_ _12364_/A _11493_/B VGND VGND VPWR VPWR _11493_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16020_ _15942_/X _16020_/B VGND VGND VPWR VPWR _16020_/Y sky130_fd_sc_hd__nand2b_1
X_13232_ _14528_/A VGND VGND VPWR VPWR _14736_/A sky130_fd_sc_hd__buf_1
X_10444_ _10444_/A VGND VGND VPWR VPWR _10444_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13163_ _15255_/A _13111_/B _13111_/Y VGND VGND VPWR VPWR _13163_/Y sky130_fd_sc_hd__o21ai_1
X_10375_ _10251_/A _10170_/B _10170_/Y VGND VGND VPWR VPWR _10376_/A sky130_fd_sc_hd__a21oi_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12114_ _12062_/X _12113_/Y _12062_/X _12113_/Y VGND VGND VPWR VPWR _12151_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13094_ _13011_/X _13093_/Y _13011_/X _13093_/Y VGND VGND VPWR VPWR _13103_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12045_ _12045_/A VGND VGND VPWR VPWR _12045_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15804_ _15672_/X _15803_/Y _15672_/X _15803_/Y VGND VGND VPWR VPWR _16207_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13996_ _13543_/X _13995_/Y _13543_/X _13995_/Y VGND VGND VPWR VPWR _13996_/X sky130_fd_sc_hd__a2bb2o_1
X_15735_ _15681_/A _15681_/B _15681_/Y VGND VGND VPWR VPWR _15735_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12947_ _12872_/Y _12945_/X _12946_/Y VGND VGND VPWR VPWR _12947_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15666_ _15777_/A _16028_/A _15664_/X _15778_/A VGND VGND VPWR VPWR _15666_/X sky130_fd_sc_hd__a31o_1
XFILLER_60_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12878_ _12855_/A _12855_/B _12855_/Y VGND VGND VPWR VPWR _12878_/Y sky130_fd_sc_hd__o21ai_1
X_14617_ _15343_/A _14657_/B VGND VGND VPWR VPWR _14617_/Y sky130_fd_sc_hd__nor2_1
X_11829_ _11797_/X _11828_/X _11797_/X _11828_/X VGND VGND VPWR VPWR _11840_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15597_ _14317_/X _15597_/B VGND VGND VPWR VPWR _15597_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14548_ _14548_/A _14517_/X VGND VGND VPWR VPWR _14548_/X sky130_fd_sc_hd__or2b_1
X_14479_ _15193_/A _14521_/B VGND VGND VPWR VPWR _14540_/A sky130_fd_sc_hd__and2_1
X_16218_ _16218_/A VGND VGND VPWR VPWR _16218_/Y sky130_fd_sc_hd__inv_2
X_16149_ _16147_/A _16148_/A _16147_/Y _16148_/Y _16388_/A VGND VGND VPWR VPWR _16270_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08971_ _08912_/X _08969_/X _11391_/B VGND VGND VPWR VPWR _08971_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09523_ _09521_/Y _09522_/X _09521_/Y _09522_/X VGND VGND VPWR VPWR _09523_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_101_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09454_ _09492_/A _09454_/B VGND VGND VPWR VPWR _09454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09385_ _09431_/B _09376_/B _09376_/X _11271_/A VGND VGND VPWR VPWR _11476_/A sky130_fd_sc_hd__a22o_1
X_08405_ _08653_/A VGND VGND VPWR VPWR _08944_/A sky130_fd_sc_hd__inv_2
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08336_ _08336_/A input31/X VGND VGND VPWR VPWR _08337_/B sky130_fd_sc_hd__nor2_1
X_08267_ input12/X VGND VGND VPWR VPWR _08352_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10160_ _10114_/A _10114_/B _10115_/A VGND VGND VPWR VPWR _10163_/A sky130_fd_sc_hd__a21bo_1
XFILLER_126_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10091_ _09194_/Y _10090_/X _09194_/Y _10090_/X VGND VGND VPWR VPWR _10091_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13850_ _13814_/Y _13848_/X _13849_/Y VGND VGND VPWR VPWR _13850_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13781_ _13781_/A VGND VGND VPWR VPWR _13781_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12801_ _12779_/X _12800_/Y _12779_/X _12800_/Y VGND VGND VPWR VPWR _12855_/B sky130_fd_sc_hd__a2bb2o_1
X_10993_ _10954_/X _10992_/X _10954_/X _10992_/X VGND VGND VPWR VPWR _11122_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15520_ _15639_/A _15640_/A _15519_/X VGND VGND VPWR VPWR _15524_/B sky130_fd_sc_hd__o21ai_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12732_ _12718_/X _12731_/X _12718_/X _12731_/X VGND VGND VPWR VPWR _12782_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15451_ _15409_/X _15450_/X _15409_/X _15450_/X VGND VGND VPWR VPWR _15452_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14402_ _15972_/A _14402_/B VGND VGND VPWR VPWR _14402_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12663_/A VGND VGND VPWR VPWR _12663_/Y sky130_fd_sc_hd__inv_2
X_12594_ _12620_/A _12620_/B VGND VGND VPWR VPWR _12594_/X sky130_fd_sc_hd__and2_1
X_15382_ _15336_/X _15381_/X _15336_/X _15381_/X VGND VGND VPWR VPWR _15404_/B sky130_fd_sc_hd__a2bb2o_1
X_11614_ _11614_/A VGND VGND VPWR VPWR _11614_/X sky130_fd_sc_hd__buf_1
XFILLER_7_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14333_ _13429_/Y _14332_/X _13429_/Y _14332_/X VGND VGND VPWR VPWR _14334_/B sky130_fd_sc_hd__a2bb2oi_1
X_11545_ _11635_/A _11544_/Y _11635_/A _11544_/Y VGND VGND VPWR VPWR _11641_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14264_ _14264_/A VGND VGND VPWR VPWR _14264_/Y sky130_fd_sc_hd__inv_2
X_11476_ _11476_/A _11476_/B VGND VGND VPWR VPWR _11476_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16003_ _15961_/X _16002_/Y _15961_/X _16002_/Y VGND VGND VPWR VPWR _16044_/B sky130_fd_sc_hd__a2bb2o_1
X_13215_ _14858_/A _13306_/B VGND VGND VPWR VPWR _13215_/Y sky130_fd_sc_hd__nor2_1
X_10427_ _12234_/A _11795_/B VGND VGND VPWR VPWR _10625_/A sky130_fd_sc_hd__nand2_1
X_14195_ _14195_/A _12630_/X VGND VGND VPWR VPWR _14195_/X sky130_fd_sc_hd__or2b_1
XFILLER_112_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13146_ _13122_/X _13145_/Y _13122_/X _13145_/Y VGND VGND VPWR VPWR _13204_/B sky130_fd_sc_hd__a2bb2o_1
X_10358_ _15028_/A _10338_/B _10338_/X _10357_/X VGND VGND VPWR VPWR _10358_/X sky130_fd_sc_hd__o22a_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13077_ _15255_/A _13111_/B VGND VGND VPWR VPWR _13077_/Y sky130_fd_sc_hd__nor2_1
X_10289_ _10289_/A _10352_/A VGND VGND VPWR VPWR _10289_/X sky130_fd_sc_hd__or2_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12028_ _13192_/A _12059_/B VGND VGND VPWR VPWR _12028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13979_ _13977_/X _13979_/B VGND VGND VPWR VPWR _13979_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_46_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15718_ _16121_/A _15819_/B VGND VGND VPWR VPWR _15718_/X sky130_fd_sc_hd__and2_1
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15649_ _15512_/A _15512_/B _15512_/X VGND VGND VPWR VPWR _15650_/A sky130_fd_sc_hd__o21ba_1
X_09170_ _09750_/A VGND VGND VPWR VPWR _09429_/A sky130_fd_sc_hd__buf_1
XFILLER_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08954_ _10018_/A _10124_/A _08836_/Y VGND VGND VPWR VPWR _08954_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08885_ _08980_/A _08980_/B VGND VGND VPWR VPWR _08885_/X sky130_fd_sc_hd__and2_1
XFILLER_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09506_ _08922_/A _09503_/Y _09503_/A _09505_/Y VGND VGND VPWR VPWR _09506_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09437_ _09322_/A _09435_/Y _09436_/Y VGND VGND VPWR VPWR _11107_/A sky130_fd_sc_hd__o21ai_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09368_ _09336_/X _08873_/Y _09336_/X _08873_/Y VGND VGND VPWR VPWR _10238_/A sky130_fd_sc_hd__o2bb2a_1
X_09299_ _09297_/A _09297_/B _09296_/Y _09298_/Y VGND VGND VPWR VPWR _09303_/A sky130_fd_sc_hd__o22a_1
X_08319_ _08319_/A VGND VGND VPWR VPWR _08319_/Y sky130_fd_sc_hd__inv_2
X_11330_ _09376_/B _10239_/B _10239_/X VGND VGND VPWR VPWR _11331_/B sky130_fd_sc_hd__a21boi_1
XFILLER_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11261_ _15449_/A _11197_/B _11197_/Y _11260_/X VGND VGND VPWR VPWR _11261_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11192_ _13364_/A VGND VGND VPWR VPWR _14017_/A sky130_fd_sc_hd__inv_2
X_13000_ _13014_/A _13015_/B VGND VGND VPWR VPWR _13090_/A sky130_fd_sc_hd__and2_1
X_10212_ _10282_/A _11724_/A _10281_/A VGND VGND VPWR VPWR _10212_/X sky130_fd_sc_hd__o21a_1
XFILLER_121_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10143_ _10143_/A _10143_/B VGND VGND VPWR VPWR _10143_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14951_ _14976_/A _14976_/B VGND VGND VPWR VPWR _14951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10074_ _10023_/X _10073_/Y _10023_/X _10073_/Y VGND VGND VPWR VPWR _10075_/B sky130_fd_sc_hd__a2bb2o_1
X_14882_ _14822_/X _14881_/X _14822_/X _14881_/X VGND VGND VPWR VPWR _14918_/B sky130_fd_sc_hd__a2bb2o_1
X_13902_ _14610_/A _13853_/B _13853_/Y VGND VGND VPWR VPWR _13902_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13833_ _13837_/A VGND VGND VPWR VPWR _14643_/A sky130_fd_sc_hd__buf_1
XFILLER_63_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15503_ _15544_/A _15544_/B VGND VGND VPWR VPWR _15503_/X sky130_fd_sc_hd__and2_1
X_13764_ _13764_/A _13764_/B VGND VGND VPWR VPWR _13764_/X sky130_fd_sc_hd__or2_1
XFILLER_71_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10976_ _10976_/A VGND VGND VPWR VPWR _11529_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13695_ _13735_/A _13693_/X _13694_/X VGND VGND VPWR VPWR _13695_/X sky130_fd_sc_hd__o21a_1
X_12715_ _12695_/A _12695_/B _12695_/Y _12714_/X VGND VGND VPWR VPWR _12715_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12646_ _15554_/A VGND VGND VPWR VPWR _14984_/A sky130_fd_sc_hd__buf_1
X_15434_ _15563_/A _15563_/B _15433_/Y VGND VGND VPWR VPWR _15434_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15365_ _15416_/A _15416_/B VGND VGND VPWR VPWR _15441_/A sky130_fd_sc_hd__and2_1
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14316_ _14270_/A _14315_/Y _14270_/A _14315_/Y VGND VGND VPWR VPWR _14391_/B sky130_fd_sc_hd__a2bb2o_1
X_12577_ _15524_/A VGND VGND VPWR VPWR _14910_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15296_ _15351_/A _15351_/B VGND VGND VPWR VPWR _15296_/X sky130_fd_sc_hd__and2_1
XFILLER_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11528_ rebuffer22/X _11527_/Y _11528_/B1 _11527_/Y VGND VGND VPWR VPWR _11529_/B
+ sky130_fd_sc_hd__a2bb2oi_1
X_14247_ _14247_/A _15838_/A VGND VGND VPWR VPWR _14248_/B sky130_fd_sc_hd__nand2_1
X_11459_ _14125_/A _11372_/B _11372_/Y _12524_/A VGND VGND VPWR VPWR _12516_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14178_ _12635_/X _14177_/X _12635_/X _14177_/X VGND VGND VPWR VPWR _14277_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13129_ _12954_/A _13036_/X _12953_/X VGND VGND VPWR VPWR _13129_/X sky130_fd_sc_hd__o21a_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08670_ _08670_/A VGND VGND VPWR VPWR _08929_/A sky130_fd_sc_hd__inv_4
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09222_ _09802_/A VGND VGND VPWR VPWR _09693_/A sky130_fd_sc_hd__inv_2
XFILLER_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09153_ _08762_/A _09147_/X _09147_/X _08535_/Y VGND VGND VPWR VPWR _09154_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_107_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09084_ _09766_/A VGND VGND VPWR VPWR _09426_/A sky130_fd_sc_hd__buf_1
XFILLER_103_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09986_ _09986_/A _09987_/B VGND VGND VPWR VPWR _09986_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08937_ _09041_/A _08937_/B VGND VGND VPWR VPWR _08937_/X sky130_fd_sc_hd__or2_1
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08868_ _09482_/A _08760_/Y _08762_/Y _08867_/X VGND VGND VPWR VPWR _08868_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08799_ _08798_/X _08731_/Y _08798_/A _08731_/Y VGND VGND VPWR VPWR _08801_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10830_ _10829_/A _10829_/B _10829_/Y _10984_/A VGND VGND VPWR VPWR _12082_/A sky130_fd_sc_hd__o211a_1
X_10761_ _10766_/A _10760_/X _10766_/A _10760_/X VGND VGND VPWR VPWR _10769_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12500_ _12649_/A VGND VGND VPWR VPWR _12501_/A sky130_fd_sc_hd__inv_2
X_13480_ _13480_/A VGND VGND VPWR VPWR _13480_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10692_ _10692_/A _10692_/B VGND VGND VPWR VPWR _10692_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12431_ _12431_/A _12435_/B VGND VGND VPWR VPWR _12431_/X sky130_fd_sc_hd__or2_1
XFILLER_126_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12362_ _13043_/A _12362_/B VGND VGND VPWR VPWR _12362_/Y sky130_fd_sc_hd__nor2_1
X_15150_ _15137_/A _15137_/B _15137_/Y _15149_/X VGND VGND VPWR VPWR _15150_/X sky130_fd_sc_hd__a2bb2o_1
X_14101_ _14097_/Y _14099_/Y _14100_/Y VGND VGND VPWR VPWR _14105_/B sky130_fd_sc_hd__o21ai_1
X_12293_ _13204_/A _12360_/B _12292_/Y VGND VGND VPWR VPWR _12293_/Y sky130_fd_sc_hd__o21ai_1
X_15081_ _15081_/A _15081_/B VGND VGND VPWR VPWR _15081_/Y sky130_fd_sc_hd__nand2_1
X_11313_ _12268_/A VGND VGND VPWR VPWR _12181_/A sky130_fd_sc_hd__inv_2
XFILLER_107_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11244_ _12232_/A _11244_/B VGND VGND VPWR VPWR _11244_/Y sky130_fd_sc_hd__nand2_1
X_14032_ _14032_/A VGND VGND VPWR VPWR _15464_/A sky130_fd_sc_hd__buf_1
XFILLER_106_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11175_ _13893_/A _11176_/B VGND VGND VPWR VPWR _11177_/A sky130_fd_sc_hd__and2_1
XFILLER_79_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15983_ _15973_/X _15981_/X _15988_/B VGND VGND VPWR VPWR _15983_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10126_ _10126_/A _10126_/B VGND VGND VPWR VPWR _10127_/B sky130_fd_sc_hd__or2_1
XFILLER_121_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14934_ _14934_/A VGND VGND VPWR VPWR _14971_/A sky130_fd_sc_hd__clkbuf_2
X_10057_ _08843_/A _09070_/A _08944_/X VGND VGND VPWR VPWR _10057_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14865_ _14774_/A _14774_/B _14774_/A _14774_/B VGND VGND VPWR VPWR _14865_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14796_ _14796_/A _14730_/X VGND VGND VPWR VPWR _14796_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13816_ _13763_/X _13815_/X _13763_/X _13815_/X VGND VGND VPWR VPWR _13847_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13747_ _14500_/A _13686_/B _13686_/Y VGND VGND VPWR VPWR _13747_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10959_ _10959_/A VGND VGND VPWR VPWR _10959_/X sky130_fd_sc_hd__clkbuf_2
X_16466_ _08229_/A _16466_/D VGND VGND VPWR VPWR _16466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15417_ _15441_/A _15415_/X _15416_/X VGND VGND VPWR VPWR _15417_/X sky130_fd_sc_hd__o21a_1
X_13678_ _13617_/X _13677_/X _13617_/X _13677_/X VGND VGND VPWR VPWR _13686_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16397_ _16397_/A _16397_/B _16397_/C _16397_/D VGND VGND VPWR VPWR _16407_/B sky130_fd_sc_hd__or4_2
X_12629_ _14201_/A _12627_/X _12628_/X VGND VGND VPWR VPWR _12629_/X sky130_fd_sc_hd__o21a_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15348_ _15366_/A _15346_/X _15347_/X VGND VGND VPWR VPWR _15348_/X sky130_fd_sc_hd__o21a_1
X_15279_ _14585_/A _15249_/B _15249_/Y _15278_/X VGND VGND VPWR VPWR _15279_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _09687_/A _09834_/Y _09801_/B VGND VGND VPWR VPWR _10499_/A sky130_fd_sc_hd__o21ai_2
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09700_/A _09770_/Y _09725_/Y VGND VGND VPWR VPWR _09773_/B sky130_fd_sc_hd__o21ai_1
XFILLER_112_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08722_ _08852_/A _09540_/A _09234_/A _09041_/A VGND VGND VPWR VPWR _08722_/X sky130_fd_sc_hd__o22a_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08653_ _08653_/A VGND VGND VPWR VPWR _08843_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _08584_/A VGND VGND VPWR VPWR _10115_/B sky130_fd_sc_hd__inv_2
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09205_ _09040_/Y _09145_/A _09040_/A _09145_/Y _09204_/X VGND VGND VPWR VPWR _13368_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09136_ _09426_/A _09136_/B VGND VGND VPWR VPWR _09136_/Y sky130_fd_sc_hd__nand2_1
X_09067_ _08930_/A _09829_/A _08922_/A VGND VGND VPWR VPWR _09627_/A sky130_fd_sc_hd__o21ai_2
XFILLER_104_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09969_ _10077_/A VGND VGND VPWR VPWR _09969_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12980_ _13696_/A VGND VGND VPWR VPWR _14480_/A sky130_fd_sc_hd__inv_2
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11931_ _12776_/A _11988_/A VGND VGND VPWR VPWR _11931_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14650_ _14633_/Y _14648_/X _14649_/Y VGND VGND VPWR VPWR _14650_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11862_ _11862_/A _11862_/B VGND VGND VPWR VPWR _11863_/B sky130_fd_sc_hd__or2_1
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14581_ _14581_/A _14581_/B VGND VGND VPWR VPWR _14581_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13601_ _13620_/A _13621_/B VGND VGND VPWR VPWR _13601_/Y sky130_fd_sc_hd__nor2_1
X_10813_ _10810_/Y _12693_/A _10676_/X _10812_/Y VGND VGND VPWR VPWR _10813_/X sky130_fd_sc_hd__o22a_1
X_16320_ _16320_/A _16320_/B VGND VGND VPWR VPWR _16320_/Y sky130_fd_sc_hd__nand2_1
X_11793_ _10426_/B _11792_/Y _10426_/B _11792_/Y VGND VGND VPWR VPWR _11794_/B sky130_fd_sc_hd__a2bb2o_1
X_13532_ _15030_/A _13527_/B _13527_/Y _13531_/X VGND VGND VPWR VPWR _13532_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10744_ _10744_/A VGND VGND VPWR VPWR _10744_/Y sky130_fd_sc_hd__inv_2
X_16251_ _16251_/A _16251_/B VGND VGND VPWR VPWR _16251_/Y sky130_fd_sc_hd__nand2_1
X_13463_ _15422_/A _12789_/B _12789_/Y _12862_/X VGND VGND VPWR VPWR _13463_/X sky130_fd_sc_hd__o2bb2a_1
X_10675_ _10675_/A _11862_/A VGND VGND VPWR VPWR _10675_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16182_ _16110_/A _15811_/B _15811_/Y VGND VGND VPWR VPWR _16182_/X sky130_fd_sc_hd__o21a_1
X_13394_ _14102_/A VGND VGND VPWR VPWR _14105_/A sky130_fd_sc_hd__buf_1
X_15202_ _15202_/A _15202_/B VGND VGND VPWR VPWR _15202_/Y sky130_fd_sc_hd__nand2_1
X_12414_ _13494_/A VGND VGND VPWR VPWR _13457_/A sky130_fd_sc_hd__buf_1
X_12345_ _12243_/X _12344_/Y _12243_/X _12344_/Y VGND VGND VPWR VPWR _12561_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15133_ _15091_/X _15132_/Y _15091_/X _15132_/Y VGND VGND VPWR VPWR _15134_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15064_ _15064_/A _15040_/X VGND VGND VPWR VPWR _15064_/X sky130_fd_sc_hd__or2b_1
X_12276_ _12274_/X _12276_/B VGND VGND VPWR VPWR _12276_/Y sky130_fd_sc_hd__nand2b_1
X_11227_ _13340_/A VGND VGND VPWR VPWR _14032_/A sky130_fd_sc_hd__inv_2
X_14015_ _15412_/A _13953_/B _13953_/Y VGND VGND VPWR VPWR _14015_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11158_ _11314_/A _12268_/A _11157_/Y VGND VGND VPWR VPWR _11158_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10109_ _10109_/A VGND VGND VPWR VPWR _10109_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15966_ _15966_/A _15966_/B VGND VGND VPWR VPWR _15966_/Y sky130_fd_sc_hd__nand2_1
X_11089_ _11211_/A _11087_/X _11088_/X VGND VGND VPWR VPWR _11089_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15897_ _15868_/Y _15895_/X _15896_/Y VGND VGND VPWR VPWR _15897_/X sky130_fd_sc_hd__o21a_1
X_14917_ _14886_/Y _14915_/X _14916_/Y VGND VGND VPWR VPWR _14917_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14848_ _15178_/A _14848_/B VGND VGND VPWR VPWR _14848_/X sky130_fd_sc_hd__or2_1
XFILLER_91_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14779_ _15446_/A VGND VGND VPWR VPWR _14782_/A sky130_fd_sc_hd__buf_1
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16449_ _16412_/Y _16473_/Q _16446_/Y _16428_/Y VGND VGND VPWR VPWR _16449_/X sky130_fd_sc_hd__o211a_1
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09823_ _09820_/A _09820_/B _09821_/B VGND VGND VPWR VPWR _09848_/A sky130_fd_sc_hd__a21bo_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09754_ _09754_/A VGND VGND VPWR VPWR _09788_/A sky130_fd_sc_hd__inv_2
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09685_ _08645_/X _09687_/B _08645_/A _09687_/B VGND VGND VPWR VPWR _09686_/B sky130_fd_sc_hd__a2bb2o_1
X_08705_ _09341_/A VGND VGND VPWR VPWR _08706_/B sky130_fd_sc_hd__inv_2
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _09462_/B _10111_/B VGND VGND VPWR VPWR _08637_/A sky130_fd_sc_hd__or2_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08567_ _09734_/A _08567_/B VGND VGND VPWR VPWR _08567_/X sky130_fd_sc_hd__or2_1
X_08498_ _08660_/A VGND VGND VPWR VPWR _08650_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10460_ _10460_/A VGND VGND VPWR VPWR _10460_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09119_ _09115_/Y _09117_/Y _09118_/Y VGND VGND VPWR VPWR _09123_/B sky130_fd_sc_hd__o21ai_1
XFILLER_129_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10391_ _10360_/X _10390_/X _10360_/X _10390_/X VGND VGND VPWR VPWR _10392_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12130_ _12141_/A _12141_/B VGND VGND VPWR VPWR _12227_/A sky130_fd_sc_hd__and2_1
X_12061_ _12061_/A _12061_/B VGND VGND VPWR VPWR _12061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11012_ _15063_/A VGND VGND VPWR VPWR _13901_/A sky130_fd_sc_hd__buf_1
XFILLER_77_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15820_ _15718_/X _15818_/X _16150_/B VGND VGND VPWR VPWR _15820_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15751_ _14913_/X _15750_/X _14913_/X _15750_/X VGND VGND VPWR VPWR _15752_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_100_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12963_ _14749_/A _13033_/B VGND VGND VPWR VPWR _13045_/A sky130_fd_sc_hd__and2_1
XFILLER_18_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15682_ _15599_/Y _15680_/X _15681_/Y VGND VGND VPWR VPWR _15682_/X sky130_fd_sc_hd__o21a_1
X_14702_ _15339_/A _14653_/B _14653_/Y VGND VGND VPWR VPWR _14702_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_85_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11914_ _13551_/A _11914_/B VGND VGND VPWR VPWR _11914_/X sky130_fd_sc_hd__and2_1
XFILLER_18_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14633_ _15335_/A _14649_/B VGND VGND VPWR VPWR _14633_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12894_ _12847_/A _12847_/B _12847_/Y VGND VGND VPWR VPWR _12894_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11845_ _11824_/Y _11843_/X _11844_/Y VGND VGND VPWR VPWR _11845_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14564_/A _14509_/X VGND VGND VPWR VPWR _14564_/X sky130_fd_sc_hd__or2b_1
X_11776_ _12768_/A _11775_/B _11775_/Y VGND VGND VPWR VPWR _11776_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16303_ _16255_/A _16322_/A _16255_/Y VGND VGND VPWR VPWR _16303_/Y sky130_fd_sc_hd__o21ai_1
X_14495_ _15205_/A _14513_/B VGND VGND VPWR VPWR _14556_/A sky130_fd_sc_hd__and2_1
X_13515_ _13515_/A _13515_/B VGND VGND VPWR VPWR _13515_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10727_ _10727_/A VGND VGND VPWR VPWR _10727_/Y sky130_fd_sc_hd__inv_2
X_16234_ _16234_/A VGND VGND VPWR VPWR _16234_/Y sky130_fd_sc_hd__clkinvlp_2
X_13446_ _13380_/Y _13444_/X _13445_/Y VGND VGND VPWR VPWR _13446_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10658_ _10656_/Y _10657_/Y _10657_/B _09907_/B _10794_/A VGND VGND VPWR VPWR _12938_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16165_ _16189_/A _16165_/B VGND VGND VPWR VPWR _16266_/A sky130_fd_sc_hd__or2_1
X_13377_ _14143_/A _13447_/B VGND VGND VPWR VPWR _13377_/Y sky130_fd_sc_hd__nor2_1
X_10589_ _10532_/X _10588_/Y _10532_/X _10588_/Y VGND VGND VPWR VPWR _10645_/B sky130_fd_sc_hd__a2bb2o_1
X_16096_ _16096_/A _16099_/B VGND VGND VPWR VPWR _16096_/Y sky130_fd_sc_hd__nor2_1
X_12328_ _12331_/A _12331_/B VGND VGND VPWR VPWR _12591_/A sky130_fd_sc_hd__and2_1
X_15116_ _15116_/A _15116_/B VGND VGND VPWR VPWR _15116_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12259_ _13715_/A _12259_/B VGND VGND VPWR VPWR _12259_/Y sky130_fd_sc_hd__nor2_1
X_15047_ _15055_/A _15045_/X _15046_/X VGND VGND VPWR VPWR _15047_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15949_ _15945_/X _15947_/Y _16023_/B VGND VGND VPWR VPWR _15949_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09470_ _09470_/A _09470_/B VGND VGND VPWR VPWR _09470_/X sky130_fd_sc_hd__or2_1
XFILLER_63_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08421_ _09217_/A VGND VGND VPWR VPWR _08715_/A sky130_fd_sc_hd__inv_2
XFILLER_24_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08352_ input28/X _08352_/B VGND VGND VPWR VPWR _08353_/B sky130_fd_sc_hd__nor2_1
X_08283_ _08276_/Y input25/X _08279_/Y _08399_/B VGND VGND VPWR VPWR _08389_/A sky130_fd_sc_hd__o22a_1
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09806_ _09855_/B VGND VGND VPWR VPWR _09806_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09737_ _09737_/A _09737_/B VGND VGND VPWR VPWR _09740_/B sky130_fd_sc_hd__or2_1
XFILLER_67_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09668_ _09569_/A _09569_/B _09569_/Y _09667_/Y VGND VGND VPWR VPWR _09668_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_91_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09599_ _09511_/X _09598_/X _09511_/X _09598_/X VGND VGND VPWR VPWR _09983_/A sky130_fd_sc_hd__a2bb2o_1
X_08619_ _08618_/X _08413_/Y _08618_/X _08413_/Y VGND VGND VPWR VPWR _08622_/A sky130_fd_sc_hd__o2bb2a_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _13495_/A _11629_/B _11629_/X _11511_/X VGND VGND VPWR VPWR _11630_/X sky130_fd_sc_hd__o22a_1
XFILLER_11_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11561_ _13544_/A _11561_/B VGND VGND VPWR VPWR _11561_/X sky130_fd_sc_hd__or2_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13300_ _14740_/A _13300_/B VGND VGND VPWR VPWR _13300_/Y sky130_fd_sc_hd__nand2_1
X_10512_ _10430_/X _10511_/X _10430_/X _10511_/X VGND VGND VPWR VPWR _10525_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14280_ _14133_/X _14279_/Y _14133_/X _14279_/Y VGND VGND VPWR VPWR _14281_/B sky130_fd_sc_hd__a2bb2oi_1
X_11492_ _12396_/A VGND VGND VPWR VPWR _13882_/A sky130_fd_sc_hd__buf_1
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13231_ _15063_/A VGND VGND VPWR VPWR _14528_/A sky130_fd_sc_hd__inv_2
X_10443_ _09978_/A _09978_/B _09978_/Y VGND VGND VPWR VPWR _10444_/A sky130_fd_sc_hd__o21ai_1
XFILLER_109_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13162_ _13194_/A _13194_/B VGND VGND VPWR VPWR _13162_/Y sky130_fd_sc_hd__nor2_1
X_10374_ _10374_/A VGND VGND VPWR VPWR _11808_/A sky130_fd_sc_hd__inv_4
XFILLER_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12113_ _13196_/A _12063_/B _12063_/Y VGND VGND VPWR VPWR _12113_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13093_ _13676_/A _13012_/B _13012_/Y VGND VGND VPWR VPWR _13093_/Y sky130_fd_sc_hd__o21ai_1
X_12044_ _12044_/A VGND VGND VPWR VPWR _12045_/A sky130_fd_sc_hd__buf_1
XFILLER_49_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15803_ _15673_/A _15673_/B _15673_/Y VGND VGND VPWR VPWR _15803_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15734_ _15752_/A _15734_/B VGND VGND VPWR VPWR _16112_/A sky130_fd_sc_hd__nor2_1
X_13995_ _13962_/X _13993_/Y _13994_/Y VGND VGND VPWR VPWR _13995_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12946_ _12946_/A _12946_/B VGND VGND VPWR VPWR _12946_/Y sky130_fd_sc_hd__nand2_1
X_15665_ _15665_/A _15665_/B VGND VGND VPWR VPWR _15778_/A sky130_fd_sc_hd__and2_1
X_12877_ _12942_/A VGND VGND VPWR VPWR _14599_/A sky130_fd_sc_hd__buf_1
XFILLER_61_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15596_ _16044_/A VGND VGND VPWR VPWR _15681_/A sky130_fd_sc_hd__inv_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14584_/X _14615_/Y _14584_/X _14615_/Y VGND VGND VPWR VPWR _14657_/B sky130_fd_sc_hd__a2bb2o_1
X_11828_ _10405_/A _11783_/B _10405_/A _11783_/B VGND VGND VPWR VPWR _11828_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _15255_/A VGND VGND VPWR VPWR _14581_/A sky130_fd_sc_hd__buf_1
XFILLER_119_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11759_ _11801_/A VGND VGND VPWR VPWR _12770_/A sky130_fd_sc_hd__buf_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14478_ _14469_/X _14477_/X _14469_/X _14477_/X VGND VGND VPWR VPWR _14521_/B sky130_fd_sc_hd__a2bb2o_1
X_16217_ _16217_/A VGND VGND VPWR VPWR _16217_/Y sky130_fd_sc_hd__inv_2
X_13429_ _13359_/X _13428_/X _13359_/X _13428_/X VGND VGND VPWR VPWR _13429_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16148_ _16148_/A VGND VGND VPWR VPWR _16148_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16079_ _16106_/A _16106_/B VGND VGND VPWR VPWR _16079_/X sky130_fd_sc_hd__and2_1
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08970_ _08970_/A _08970_/B VGND VGND VPWR VPWR _11391_/B sky130_fd_sc_hd__or2_1
XFILLER_102_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 wb_rst_i VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09522_ _09937_/A _09199_/Y _08703_/A _09199_/A VGND VGND VPWR VPWR _09522_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09453_ _09490_/A _09453_/B VGND VGND VPWR VPWR _09453_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09384_ _09432_/B _09382_/B _09382_/X _11097_/A VGND VGND VPWR VPWR _11271_/A sky130_fd_sc_hd__a22o_1
X_08404_ _08361_/Y _08388_/Y _08361_/A _08388_/A _08419_/A VGND VGND VPWR VPWR _08653_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08335_ _08333_/Y _08334_/A _08333_/A _08334_/Y _08304_/A VGND VGND VPWR VPWR _09209_/B
+ sky130_fd_sc_hd__o221a_1
X_08266_ _08266_/A input13/X VGND VGND VPWR VPWR _08347_/A sky130_fd_sc_hd__nor2_1
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10090_ _10031_/X _10089_/X _10031_/X _10089_/X VGND VGND VPWR VPWR _10090_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12800_ _12780_/A _12780_/B _12780_/Y VGND VGND VPWR VPWR _12800_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13780_ _13780_/A VGND VGND VPWR VPWR _15113_/A sky130_fd_sc_hd__buf_1
X_10992_ _09395_/A _11128_/B _09395_/A _11128_/B VGND VGND VPWR VPWR _10992_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _12687_/A _12687_/B _12687_/Y VGND VGND VPWR VPWR _12731_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15450_ _15450_/A _15410_/X VGND VGND VPWR VPWR _15450_/X sky130_fd_sc_hd__or2b_1
XFILLER_70_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _10452_/Y _12661_/Y _10379_/Y VGND VGND VPWR VPWR _12663_/A sky130_fd_sc_hd__o21ai_1
X_14401_ _14397_/X _14399_/Y _15687_/B VGND VGND VPWR VPWR _14401_/X sky130_fd_sc_hd__o21a_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11612_/A _12426_/B _11612_/Y VGND VGND VPWR VPWR _11614_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12593_ _12590_/Y _12592_/Y _12590_/A _12592_/A _12502_/A VGND VGND VPWR VPWR _12620_/B
+ sky130_fd_sc_hd__o221a_1
X_15381_ _15381_/A _15337_/X VGND VGND VPWR VPWR _15381_/X sky130_fd_sc_hd__or2b_1
X_14332_ _14105_/A _13430_/B _13430_/Y VGND VGND VPWR VPWR _14332_/X sky130_fd_sc_hd__o21a_1
X_11544_ _13871_/A _11634_/B _11543_/Y VGND VGND VPWR VPWR _11544_/Y sky130_fd_sc_hd__o21ai_1
X_14263_ _14209_/Y _14261_/Y _14262_/Y VGND VGND VPWR VPWR _14264_/A sky130_fd_sc_hd__o21ai_2
X_11475_ _09430_/B _09370_/B _09370_/X VGND VGND VPWR VPWR _11476_/B sky130_fd_sc_hd__a21boi_1
X_16002_ _15924_/X _16002_/B VGND VGND VPWR VPWR _16002_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_109_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13214_ _13205_/X _13213_/Y _13205_/X _13213_/Y VGND VGND VPWR VPWR _13306_/B sky130_fd_sc_hd__a2bb2o_1
X_10426_ _10426_/A _10426_/B VGND VGND VPWR VPWR _11795_/B sky130_fd_sc_hd__or2_1
X_14194_ _14206_/A _14194_/B VGND VGND VPWR VPWR _15863_/A sky130_fd_sc_hd__or2_1
XFILLER_112_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13145_ _15237_/A _13123_/B _13123_/Y VGND VGND VPWR VPWR _13145_/Y sky130_fd_sc_hd__o21ai_1
X_10357_ _12832_/A _10355_/B _10354_/X _10356_/Y VGND VGND VPWR VPWR _10357_/X sky130_fd_sc_hd__o22a_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13076_ _13020_/X _13075_/X _13020_/X _13075_/X VGND VGND VPWR VPWR _13111_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _12606_/A _10288_/B VGND VGND VPWR VPWR _10352_/A sky130_fd_sc_hd__or2_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12027_ _11973_/X _12026_/Y _11973_/X _12026_/Y VGND VGND VPWR VPWR _12059_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13978_ _13978_/A _13978_/B VGND VGND VPWR VPWR _13979_/B sky130_fd_sc_hd__or2_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15717_ _15693_/Y _15716_/Y _15693_/Y _15716_/Y VGND VGND VPWR VPWR _15819_/B sky130_fd_sc_hd__a2bb2o_1
X_12929_ _12908_/Y _12927_/X _12928_/Y VGND VGND VPWR VPWR _12929_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15648_ _14376_/X _15647_/Y _14376_/X _15647_/Y VGND VGND VPWR VPWR _15667_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15579_ _15497_/X _15579_/B VGND VGND VPWR VPWR _15579_/X sky130_fd_sc_hd__and2b_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08953_ _08948_/Y _08951_/Y _08952_/Y VGND VGND VPWR VPWR _08960_/A sky130_fd_sc_hd__o21ai_1
XFILLER_69_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08884_ _08883_/Y _08865_/X _08883_/Y _08865_/X VGND VGND VPWR VPWR _08980_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09505_ _09505_/A VGND VGND VPWR VPWR _09505_/Y sky130_fd_sc_hd__inv_4
XFILLER_112_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09436_/B VGND VGND VPWR VPWR _09436_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A VGND VGND VPWR VPWR _09430_/B sky130_fd_sc_hd__inv_2
X_09298_ _09298_/A VGND VGND VPWR VPWR _09298_/Y sky130_fd_sc_hd__inv_2
X_08318_ _08318_/A VGND VGND VPWR VPWR _08318_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08249_ input3/X VGND VGND VPWR VPWR _08321_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_125_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11260_ _15452_/A _11206_/B _11206_/Y _11259_/X VGND VGND VPWR VPWR _11260_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10211_ _10462_/A _11714_/A VGND VGND VPWR VPWR _10281_/A sky130_fd_sc_hd__nand2_1
X_11191_ _09135_/Y _11190_/A _09135_/A _11190_/Y _09204_/X VGND VGND VPWR VPWR _13364_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_106_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10142_ _10132_/A _10132_/B _10133_/B VGND VGND VPWR VPWR _10143_/B sky130_fd_sc_hd__a21bo_1
X_14950_ _14935_/X _14949_/X _14935_/X _14949_/X VGND VGND VPWR VPWR _14976_/B sky130_fd_sc_hd__a2bb2o_1
X_10073_ _10073_/A _10073_/B VGND VGND VPWR VPWR _10073_/Y sky130_fd_sc_hd__nor2_1
X_14881_ _14790_/A _14790_/B _14790_/A _14790_/B VGND VGND VPWR VPWR _14881_/X sky130_fd_sc_hd__a2bb2o_1
X_13901_ _13901_/A VGND VGND VPWR VPWR _15412_/A sky130_fd_sc_hd__buf_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13832_ _13832_/A VGND VGND VPWR VPWR _13837_/A sky130_fd_sc_hd__inv_2
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13763_ _13818_/A _13761_/X _13762_/X VGND VGND VPWR VPWR _13763_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15502_ _15481_/X _15501_/X _15481_/X _15501_/X VGND VGND VPWR VPWR _15544_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12714_ _12697_/A _12697_/B _12697_/Y _12713_/X VGND VGND VPWR VPWR _12714_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10975_ _10975_/A VGND VGND VPWR VPWR _10975_/Y sky130_fd_sc_hd__inv_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13694_ _13694_/A _13694_/B VGND VGND VPWR VPWR _13694_/X sky130_fd_sc_hd__or2_1
XFILLER_31_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12645_ _12644_/A _12644_/B _12644_/Y _11710_/X VGND VGND VPWR VPWR _12651_/A sky130_fd_sc_hd__o211ai_1
X_15433_ _15433_/A _15563_/B VGND VGND VPWR VPWR _15433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12576_ _12576_/A VGND VGND VPWR VPWR _12576_/Y sky130_fd_sc_hd__inv_2
X_15364_ _15348_/X _15363_/X _15348_/X _15363_/X VGND VGND VPWR VPWR _15416_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14315_ _15860_/A _14271_/B _14271_/Y VGND VGND VPWR VPWR _14315_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11527_ _10238_/B _10139_/B _10139_/Y VGND VGND VPWR VPWR _11527_/Y sky130_fd_sc_hd__a21oi_1
X_15295_ _15282_/X _15294_/Y _15282_/X _15294_/Y VGND VGND VPWR VPWR _15351_/B sky130_fd_sc_hd__a2bb2o_1
X_14246_ _11709_/A _14361_/B _12502_/A _15781_/A VGND VGND VPWR VPWR _15838_/A sky130_fd_sc_hd__o22a_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11458_ _14119_/A _11379_/B _11379_/Y _12532_/A VGND VGND VPWR VPWR _12524_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14177_ _14177_/A _12636_/X VGND VGND VPWR VPWR _14177_/X sky130_fd_sc_hd__or2b_1
X_11389_ _11393_/A _11389_/B VGND VGND VPWR VPWR _14107_/A sky130_fd_sc_hd__or2_1
X_10409_ _11783_/A _10409_/B VGND VGND VPWR VPWR _10409_/X sky130_fd_sc_hd__and2_1
XFILLER_125_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13128_ _13038_/Y _13126_/X _13127_/Y VGND VGND VPWR VPWR _13128_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13059_ _13770_/A VGND VGND VPWR VPWR _15246_/A sky130_fd_sc_hd__buf_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09221_ _09221_/A _09221_/B VGND VGND VPWR VPWR _09802_/A sky130_fd_sc_hd__or2_1
X_09152_ _09152_/A VGND VGND VPWR VPWR _09525_/B sky130_fd_sc_hd__inv_2
XFILLER_108_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09083_ _10013_/B _09076_/B _09077_/B VGND VGND VPWR VPWR _09766_/A sky130_fd_sc_hd__a21bo_1
XFILLER_131_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09985_ _09969_/Y _09983_/Y _09984_/Y VGND VGND VPWR VPWR _09987_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08936_ _09503_/A _10103_/A _08935_/X VGND VGND VPWR VPWR _08936_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08867_ _09484_/A _08768_/Y _08770_/Y _08866_/X VGND VGND VPWR VPWR _08867_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08798_ _08798_/A VGND VGND VPWR VPWR _08798_/X sky130_fd_sc_hd__buf_1
X_10760_ _13004_/A _10629_/B _10629_/Y VGND VGND VPWR VPWR _10760_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10691_ _09268_/B _10243_/B _10243_/X VGND VGND VPWR VPWR _10692_/B sky130_fd_sc_hd__a21boi_1
X_09419_ _10437_/A _09417_/Y _09418_/Y VGND VGND VPWR VPWR _09421_/B sky130_fd_sc_hd__o21ai_1
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12430_ _12427_/X _12429_/X _12427_/X _12429_/X VGND VGND VPWR VPWR _12432_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14100_ _14100_/A _14100_/B VGND VGND VPWR VPWR _14100_/Y sky130_fd_sc_hd__nand2_1
X_12361_ _12360_/Y _12252_/X _12292_/Y VGND VGND VPWR VPWR _12361_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12292_ _12292_/A _12360_/B VGND VGND VPWR VPWR _12292_/Y sky130_fd_sc_hd__nand2_1
X_15080_ _15029_/X _15079_/X _15029_/X _15079_/X VGND VGND VPWR VPWR _15081_/B sky130_fd_sc_hd__a2bb2o_1
X_11312_ _12268_/A VGND VGND VPWR VPWR _12687_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11243_ _11076_/X _11242_/X _11076_/X _11242_/X VGND VGND VPWR VPWR _11244_/B sky130_fd_sc_hd__a2bb2o_1
X_14031_ _14031_/A _14031_/B VGND VGND VPWR VPWR _14031_/X sky130_fd_sc_hd__and2_1
XFILLER_134_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11174_ _11104_/X _11173_/X _11104_/X _11173_/X VGND VGND VPWR VPWR _11176_/B sky130_fd_sc_hd__a2bb2o_1
X_15982_ _15982_/A _15982_/B VGND VGND VPWR VPWR _15988_/B sky130_fd_sc_hd__or2_1
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10125_ _10125_/A _10125_/B VGND VGND VPWR VPWR _10126_/B sky130_fd_sc_hd__or2_1
XFILLER_121_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14933_ _14829_/X _14859_/A _14858_/X VGND VGND VPWR VPWR _14933_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10056_ _10055_/A _10055_/B _09954_/Y _10055_/X VGND VGND VPWR VPWR _10059_/A sky130_fd_sc_hd__a22o_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14864_ _14864_/A VGND VGND VPWR VPWR _15550_/A sky130_fd_sc_hd__buf_1
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14795_ _15458_/A VGND VGND VPWR VPWR _14798_/A sky130_fd_sc_hd__buf_1
X_13815_ _13815_/A _13764_/X VGND VGND VPWR VPWR _13815_/X sky130_fd_sc_hd__or2b_1
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13746_ _13758_/A _13758_/B VGND VGND VPWR VPWR _13825_/A sky130_fd_sc_hd__and2_1
XFILLER_44_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10958_ _10958_/A VGND VGND VPWR VPWR _10958_/Y sky130_fd_sc_hd__inv_2
X_16465_ _16357_/A _16465_/D VGND VGND VPWR VPWR _16465_/Q sky130_fd_sc_hd__dfxtp_1
X_13677_ _12925_/A _13608_/B _12925_/A _13608_/B VGND VGND VPWR VPWR _13677_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12628_ _12628_/A _12628_/B VGND VGND VPWR VPWR _12628_/X sky130_fd_sc_hd__or2_1
X_15416_ _15416_/A _15416_/B VGND VGND VPWR VPWR _15416_/X sky130_fd_sc_hd__or2_1
X_10889_ _10402_/A _10888_/Y _10402_/Y _10888_/A _09445_/A VGND VGND VPWR VPWR _12053_/A
+ sky130_fd_sc_hd__a221o_2
X_16396_ _16396_/A _16396_/B _16396_/C _16457_/S VGND VGND VPWR VPWR _16397_/B sky130_fd_sc_hd__or4b_1
XFILLER_8_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12559_ _12559_/A VGND VGND VPWR VPWR _12559_/Y sky130_fd_sc_hd__inv_2
X_15347_ _15347_/A _15347_/B VGND VGND VPWR VPWR _15347_/X sky130_fd_sc_hd__or2_1
XFILLER_8_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15278_ _14583_/A _15252_/B _15252_/Y _15277_/X VGND VGND VPWR VPWR _15278_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14229_ _14085_/Y _14228_/X _14085_/Y _14228_/X VGND VGND VPWR VPWR _14230_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_7_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09770_/A _09770_/B VGND VGND VPWR VPWR _09770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08721_/A _08721_/B VGND VGND VPWR VPWR _09041_/A sky130_fd_sc_hd__nor2_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08652_ _08721_/B VGND VGND VPWR VPWR _08679_/A sky130_fd_sc_hd__buf_1
XFILLER_66_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08583_ _08714_/B VGND VGND VPWR VPWR _09467_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09204_ _11220_/B VGND VGND VPWR VPWR _09204_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09135_ _09135_/A VGND VGND VPWR VPWR _09135_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09066_ _09066_/A VGND VGND VPWR VPWR _09829_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09968_ _10079_/A VGND VGND VPWR VPWR _09968_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08919_ _08919_/A VGND VGND VPWR VPWR _09541_/A sky130_fd_sc_hd__inv_2
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11930_ _11992_/B _11929_/Y _11992_/B _11929_/Y VGND VGND VPWR VPWR _11988_/A sky130_fd_sc_hd__a2bb2o_1
X_09899_ _09728_/A _09804_/Y _09857_/B VGND VGND VPWR VPWR _09899_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11861_ _11862_/A _11862_/B VGND VGND VPWR VPWR _11861_/X sky130_fd_sc_hd__and2_1
X_14580_ _14554_/Y _14578_/X _14579_/Y VGND VGND VPWR VPWR _14580_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13600_ _13575_/X _13599_/Y _13575_/X _13599_/Y VGND VGND VPWR VPWR _13621_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11792_ _12830_/A _11720_/B _11720_/Y VGND VGND VPWR VPWR _11792_/Y sky130_fd_sc_hd__a21oi_1
X_10812_ _10812_/A _11928_/A VGND VGND VPWR VPWR _10812_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13531_ _15028_/A _13529_/B _13529_/Y _13530_/X VGND VGND VPWR VPWR _13531_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10743_ _10743_/A VGND VGND VPWR VPWR _10743_/Y sky130_fd_sc_hd__inv_2
X_16250_ _16240_/Y _16248_/Y _16249_/Y VGND VGND VPWR VPWR _16250_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13462_ _13462_/A VGND VGND VPWR VPWR _15422_/A sky130_fd_sc_hd__clkbuf_2
X_15201_ _15150_/X _15200_/Y _15150_/X _15200_/Y VGND VGND VPWR VPWR _15202_/B sky130_fd_sc_hd__a2bb2o_1
X_10674_ _11921_/A VGND VGND VPWR VPWR _11862_/A sky130_fd_sc_hd__inv_2
XFILLER_41_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16181_ _16189_/A _16181_/B VGND VGND VPWR VPWR _16262_/A sky130_fd_sc_hd__or2_1
X_13393_ _14107_/A VGND VGND VPWR VPWR _14111_/A sky130_fd_sc_hd__buf_1
X_12413_ _12413_/A VGND VGND VPWR VPWR _13494_/A sky130_fd_sc_hd__clkbuf_2
X_12344_ _12220_/A _12220_/B _12220_/Y VGND VGND VPWR VPWR _12344_/Y sky130_fd_sc_hd__o21ai_1
X_15132_ _15075_/A _15075_/B _15075_/Y VGND VGND VPWR VPWR _15132_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15063_ _15063_/A _15063_/B VGND VGND VPWR VPWR _15063_/Y sky130_fd_sc_hd__nand2_1
X_14014_ _14014_/A _14059_/B VGND VGND VPWR VPWR _14122_/A sky130_fd_sc_hd__and2_1
X_12275_ _12275_/A _12275_/B VGND VGND VPWR VPWR _12276_/B sky130_fd_sc_hd__or2_1
XFILLER_5_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11226_ _11226_/A _11251_/B VGND VGND VPWR VPWR _13340_/A sky130_fd_sc_hd__or2_1
XFILLER_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11157_ _11314_/A _12268_/A VGND VGND VPWR VPWR _11157_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10108_ _10108_/A VGND VGND VPWR VPWR _10108_/Y sky130_fd_sc_hd__clkinvlp_2
X_15965_ _15921_/X _15963_/X _15999_/B VGND VGND VPWR VPWR _15966_/B sky130_fd_sc_hd__o21a_1
X_11088_ _13909_/A _11088_/B VGND VGND VPWR VPWR _11088_/X sky130_fd_sc_hd__or2_1
XFILLER_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15896_ _15896_/A _15896_/B VGND VGND VPWR VPWR _15896_/Y sky130_fd_sc_hd__nand2_1
X_14916_ _14916_/A _14916_/B VGND VGND VPWR VPWR _14916_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10039_ _10028_/X _10038_/Y _10028_/X _10038_/Y VGND VGND VPWR VPWR _10085_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14847_ _15178_/A _14848_/B VGND VGND VPWR VPWR _14849_/A sky130_fd_sc_hd__and2_1
XFILLER_17_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14778_ _14778_/A _14778_/B VGND VGND VPWR VPWR _14778_/X sky130_fd_sc_hd__and2_1
XFILLER_51_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13729_ _13729_/A _13698_/X VGND VGND VPWR VPWR _13729_/X sky130_fd_sc_hd__or2b_1
XFILLER_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16448_ _16446_/Y _16415_/X _16412_/Y _16429_/B _16447_/X VGND VGND VPWR VPWR _16448_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16379_ _16317_/X _16378_/Y _16317_/X _16378_/Y VGND VGND VPWR VPWR _16396_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09822_ _09821_/A _09821_/B _09882_/B VGND VGND VPWR VPWR _09853_/A sky130_fd_sc_hd__a21bo_1
XFILLER_113_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09753_ _09997_/B VGND VGND VPWR VPWR _09753_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ _09937_/A _08704_/B VGND VGND VPWR VPWR _09341_/A sky130_fd_sc_hd__or2_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09684_ _09684_/A _09684_/B VGND VGND VPWR VPWR _09687_/B sky130_fd_sc_hd__or2_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08635_ _08635_/A VGND VGND VPWR VPWR _10111_/B sky130_fd_sc_hd__inv_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08566_ _09858_/A VGND VGND VPWR VPWR _09734_/A sky130_fd_sc_hd__inv_2
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08497_ _08298_/X _08496_/X _08298_/X _08496_/X VGND VGND VPWR VPWR _08660_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09118_ _09705_/A _09118_/B VGND VGND VPWR VPWR _09118_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10390_ _13521_/A _10441_/B _11758_/A _10441_/B VGND VGND VPWR VPWR _10390_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09049_ _08713_/A _08713_/B _08713_/X _09048_/Y VGND VGND VPWR VPWR _09050_/A sky130_fd_sc_hd__a22o_1
XFILLER_104_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12060_ _12028_/Y _12058_/X _12059_/Y VGND VGND VPWR VPWR _12060_/X sky130_fd_sc_hd__o21a_1
X_11011_ _12853_/A VGND VGND VPWR VPWR _15063_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15750_ _14914_/A _14914_/B _14914_/Y VGND VGND VPWR VPWR _15750_/X sky130_fd_sc_hd__o21a_1
X_12962_ _12945_/X _12961_/Y _12945_/X _12961_/Y VGND VGND VPWR VPWR _13033_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15681_ _15681_/A _15681_/B VGND VGND VPWR VPWR _15681_/Y sky130_fd_sc_hd__nand2_1
X_14701_ _14732_/A _14732_/B VGND VGND VPWR VPWR _14792_/A sky130_fd_sc_hd__and2_1
X_12893_ _12934_/A VGND VGND VPWR VPWR _14466_/A sky130_fd_sc_hd__buf_1
X_11913_ _11912_/Y _11847_/X _11870_/Y VGND VGND VPWR VPWR _11913_/X sky130_fd_sc_hd__o21a_1
X_14632_ _14576_/X _14631_/Y _14576_/X _14631_/Y VGND VGND VPWR VPWR _14649_/B sky130_fd_sc_hd__a2bb2o_1
X_11844_ _11844_/A _11844_/B VGND VGND VPWR VPWR _11844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14563_/A VGND VGND VPWR VPWR _15272_/A sky130_fd_sc_hd__buf_1
XFILLER_54_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11775_ _12768_/A _11775_/B VGND VGND VPWR VPWR _11775_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16302_ _16324_/A _16324_/B VGND VGND VPWR VPWR _16302_/Y sky130_fd_sc_hd__nor2_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14494_ _14461_/X _14493_/Y _14461_/X _14493_/Y VGND VGND VPWR VPWR _14513_/B sky130_fd_sc_hd__a2bb2o_1
X_13514_ _10575_/X _13485_/X _10575_/X _13485_/X VGND VGND VPWR VPWR _13515_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10726_ _10726_/A VGND VGND VPWR VPWR _10726_/Y sky130_fd_sc_hd__inv_2
X_16233_ _16233_/A VGND VGND VPWR VPWR _16233_/Y sky130_fd_sc_hd__clkinvlp_2
X_13445_ _13445_/A _13445_/B VGND VGND VPWR VPWR _13445_/Y sky130_fd_sc_hd__nand2_1
X_10657_ _10657_/A _10657_/B VGND VGND VPWR VPWR _10657_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16164_ _16111_/X _16163_/X _16111_/X _16163_/X VGND VGND VPWR VPWR _16165_/B sky130_fd_sc_hd__a2bb2oi_1
X_13376_ _13371_/X _13375_/X _13371_/X _13375_/X VGND VGND VPWR VPWR _13447_/B sky130_fd_sc_hd__a2bb2o_1
X_10588_ _13628_/A _10533_/B _10533_/Y VGND VGND VPWR VPWR _10588_/Y sky130_fd_sc_hd__o21ai_1
X_16095_ _16091_/Y _16213_/A _16094_/Y VGND VGND VPWR VPWR _16099_/B sky130_fd_sc_hd__o21ai_1
XFILLER_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12327_ _15512_/A _12324_/B _12324_/X _12601_/A VGND VGND VPWR VPWR _12331_/B sky130_fd_sc_hd__o22a_1
X_15115_ _15097_/X _15114_/Y _15097_/X _15114_/Y VGND VGND VPWR VPWR _15116_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12258_ _12256_/Y _12257_/Y _12192_/Y VGND VGND VPWR VPWR _12365_/A sky130_fd_sc_hd__o21ai_1
X_15046_ _15046_/A _15046_/B VGND VGND VPWR VPWR _15046_/X sky130_fd_sc_hd__or2_1
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11209_ _12217_/A VGND VGND VPWR VPWR _14023_/A sky130_fd_sc_hd__buf_1
X_12189_ _12189_/A _12259_/B VGND VGND VPWR VPWR _12189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15948_ _15948_/A _15948_/B VGND VGND VPWR VPWR _16023_/B sky130_fd_sc_hd__or2_1
XFILLER_110_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15879_ _14225_/Y _15841_/X _14225_/Y _15841_/X VGND VGND VPWR VPWR _15888_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08420_ _08418_/A _08343_/Y _08418_/Y _08343_/A _08441_/A VGND VGND VPWR VPWR _09217_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08351_ _09221_/B VGND VGND VPWR VPWR _08351_/Y sky130_fd_sc_hd__inv_2
X_08282_ _08282_/A VGND VGND VPWR VPWR _08399_/B sky130_fd_sc_hd__inv_4
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09805_ _09803_/A _09803_/B _09804_/Y VGND VGND VPWR VPWR _09855_/B sky130_fd_sc_hd__a21oi_1
XFILLER_101_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09736_ _09736_/A _09736_/B VGND VGND VPWR VPWR _09739_/A sky130_fd_sc_hd__or2_1
XFILLER_55_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09667_ _09574_/Y _09665_/X _09666_/Y VGND VGND VPWR VPWR _09667_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08618_ _09456_/A _09221_/B _10016_/A _08351_/Y VGND VGND VPWR VPWR _08618_/X sky130_fd_sc_hd__o22a_1
XFILLER_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _08795_/X _09492_/B _09492_/Y VGND VGND VPWR VPWR _09598_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08549_/A VGND VGND VPWR VPWR _08549_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_30_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11560_ _13544_/A _11561_/B VGND VGND VPWR VPWR _11562_/A sky130_fd_sc_hd__and2_1
XFILLER_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10511_ _10511_/A _10431_/X VGND VGND VPWR VPWR _10511_/X sky130_fd_sc_hd__or2b_1
XFILLER_11_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13230_ _14738_/A _13297_/B VGND VGND VPWR VPWR _13230_/Y sky130_fd_sc_hd__nor2_1
X_11491_ _11590_/A _11491_/B VGND VGND VPWR VPWR _12396_/A sky130_fd_sc_hd__nor2_2
XFILLER_108_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10442_ _13521_/A _10441_/B _10441_/X _10360_/X VGND VGND VPWR VPWR _10442_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13161_ _13112_/X _13160_/Y _13112_/X _13160_/Y VGND VGND VPWR VPWR _13194_/B sky130_fd_sc_hd__a2bb2o_1
X_10373_ _10454_/A _11220_/A VGND VGND VPWR VPWR _10374_/A sky130_fd_sc_hd__or2_1
XFILLER_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12112_ _13901_/A _12153_/B VGND VGND VPWR VPWR _12209_/A sky130_fd_sc_hd__and2_1
X_13092_ _15264_/A _13105_/B VGND VGND VPWR VPWR _13092_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12043_ _12043_/A _12043_/B VGND VGND VPWR VPWR _12044_/A sky130_fd_sc_hd__or2_1
XFILLER_104_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15802_ _16104_/A _15805_/B VGND VGND VPWR VPWR _15802_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15733_ _14919_/X _15732_/X _14919_/X _15732_/X VGND VGND VPWR VPWR _15734_/B sky130_fd_sc_hd__a2bb2oi_1
X_13994_ _13994_/A _13994_/B VGND VGND VPWR VPWR _13994_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12945_ _12876_/Y _12943_/X _12944_/Y VGND VGND VPWR VPWR _12945_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15664_ _15665_/A _15665_/B VGND VGND VPWR VPWR _15664_/X sky130_fd_sc_hd__or2_1
X_12876_ _14676_/A _12944_/B VGND VGND VPWR VPWR _12876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15595_ _15595_/A _15595_/B VGND VGND VPWR VPWR _16044_/A sky130_fd_sc_hd__or2_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _14585_/A _14585_/B _14585_/Y VGND VGND VPWR VPWR _14615_/Y sky130_fd_sc_hd__o21ai_1
X_11827_ _13620_/A _11842_/B VGND VGND VPWR VPWR _11827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _14583_/A _14583_/B VGND VGND VPWR VPWR _14546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11758_ _11758_/A VGND VGND VPWR VPWR _11801_/A sky130_fd_sc_hd__inv_2
XFILLER_14_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10709_ _09981_/A _09654_/B _09654_/Y VGND VGND VPWR VPWR _10709_/X sky130_fd_sc_hd__o21a_1
X_11689_ _11662_/A _11688_/Y _11661_/X VGND VGND VPWR VPWR _11689_/X sky130_fd_sc_hd__o21a_1
X_14477_ _14476_/A _14476_/B _14476_/Y VGND VGND VPWR VPWR _14477_/X sky130_fd_sc_hd__a21o_1
X_16216_ _16099_/A _15800_/B _15800_/Y VGND VGND VPWR VPWR _16218_/A sky130_fd_sc_hd__o21ai_1
X_13428_ _13334_/A _13334_/B _13334_/A _13334_/B VGND VGND VPWR VPWR _13428_/X sky130_fd_sc_hd__a2bb2o_1
X_16147_ _16147_/A VGND VGND VPWR VPWR _16147_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13359_ _13337_/A _13337_/B _13337_/X _13358_/X VGND VGND VPWR VPWR _13359_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16078_ _16037_/X _16077_/Y _16037_/X _16077_/Y VGND VGND VPWR VPWR _16106_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15029_ _15082_/A _15027_/X _15028_/X VGND VGND VPWR VPWR _15029_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput2 wbs_adr_i[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09521_ _09519_/Y _09520_/X _09519_/Y _09520_/X VGND VGND VPWR VPWR _09521_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_37_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09452_ _09452_/A _09531_/A VGND VGND VPWR VPWR _09452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09383_ _09327_/A _09327_/B _09327_/X _09329_/A VGND VGND VPWR VPWR _11097_/A sky130_fd_sc_hd__a22o_1
X_08403_ _08852_/A _08398_/Y _08402_/X VGND VGND VPWR VPWR _08403_/Y sky130_fd_sc_hd__o21ai_1
X_08334_ _08334_/A VGND VGND VPWR VPWR _08334_/Y sky130_fd_sc_hd__inv_2
X_08265_ input29/X VGND VGND VPWR VPWR _08266_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10991_ _10956_/X _10990_/X _10956_/X _10990_/X VGND VGND VPWR VPWR _11128_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09719_ _09720_/A _09720_/B VGND VGND VPWR VPWR _09719_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12730_ _12784_/A _12784_/B VGND VGND VPWR VPWR _12730_/Y sky130_fd_sc_hd__nor2_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12661_/A VGND VGND VPWR VPWR _12661_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14400_ _15970_/A _14400_/B VGND VGND VPWR VPWR _15687_/B sky130_fd_sc_hd__or2_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11612_/A _12426_/B VGND VGND VPWR VPWR _11612_/Y sky130_fd_sc_hd__nor2_1
X_12592_ _12592_/A VGND VGND VPWR VPWR _12592_/Y sky130_fd_sc_hd__inv_2
X_15380_ _15406_/A _15406_/B VGND VGND VPWR VPWR _15456_/A sky130_fd_sc_hd__and2_1
XFILLER_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14331_ _14261_/A _14330_/Y _14261_/A _14330_/Y VGND VGND VPWR VPWR _14385_/A sky130_fd_sc_hd__a2bb2o_1
X_11543_ _12442_/A _11634_/B VGND VGND VPWR VPWR _11543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14262_ _15869_/A _14262_/B VGND VGND VPWR VPWR _14262_/Y sky130_fd_sc_hd__nand2_1
X_11474_ _11353_/A _11269_/X _11352_/X VGND VGND VPWR VPWR _11474_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16001_ _16046_/A _16046_/B VGND VGND VPWR VPWR _16001_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14193_ _14112_/X _14192_/Y _14112_/X _14192_/Y VGND VGND VPWR VPWR _14194_/B sky130_fd_sc_hd__a2bb2oi_1
X_13213_ _13206_/A _13206_/B _13206_/Y VGND VGND VPWR VPWR _13213_/Y sky130_fd_sc_hd__o21ai_1
X_10425_ _10425_/A VGND VGND VPWR VPWR _10426_/B sky130_fd_sc_hd__inv_2
XFILLER_124_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13144_ _13206_/A _13206_/B VGND VGND VPWR VPWR _13144_/Y sky130_fd_sc_hd__nor2_1
X_10356_ _10356_/A VGND VGND VPWR VPWR _10356_/Y sky130_fd_sc_hd__inv_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13075_ _13075_/A _13021_/X VGND VGND VPWR VPWR _13075_/X sky130_fd_sc_hd__or2b_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _10287_/A VGND VGND VPWR VPWR _12606_/A sky130_fd_sc_hd__buf_2
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12026_ _11974_/A _11974_/B _11974_/Y VGND VGND VPWR VPWR _12026_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13977_ _13978_/A _13978_/B VGND VGND VPWR VPWR _13977_/X sky130_fd_sc_hd__and2_1
X_15716_ _15694_/A _15694_/B _15694_/Y VGND VGND VPWR VPWR _15716_/Y sky130_fd_sc_hd__o21ai_1
X_12928_ _12928_/A _12928_/B VGND VGND VPWR VPWR _12928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15647_ _14377_/A _14377_/B _14377_/Y VGND VGND VPWR VPWR _15647_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12859_ _12859_/A _12859_/B VGND VGND VPWR VPWR _12859_/Y sky130_fd_sc_hd__nand2_1
X_15578_ _16055_/A _15696_/B VGND VGND VPWR VPWR _15578_/Y sky130_fd_sc_hd__nor2_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14529_ _14528_/A _14528_/B _14528_/Y VGND VGND VPWR VPWR _14529_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08952_ _08952_/A _08952_/B VGND VGND VPWR VPWR _08952_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08883_ _08778_/A _10131_/A _08778_/Y VGND VGND VPWR VPWR _08883_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09504_ _08847_/A _09460_/A _09826_/B _09460_/Y VGND VGND VPWR VPWR _09505_/A sky130_fd_sc_hd__o22a_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09435_ _09763_/A _09436_/B VGND VGND VPWR VPWR _09435_/Y sky130_fd_sc_hd__nor2_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09366_ _09356_/X _09365_/X _09356_/X _09365_/X VGND VGND VPWR VPWR _09367_/A sky130_fd_sc_hd__a2bb2o_1
X_09297_ _09297_/A _09297_/B VGND VGND VPWR VPWR _09298_/A sky130_fd_sc_hd__nand2_1
X_08317_ _08317_/A _08317_/B VGND VGND VPWR VPWR _08318_/A sky130_fd_sc_hd__or2_1
X_08248_ input4/X _08248_/B VGND VGND VPWR VPWR _08317_/A sky130_fd_sc_hd__nor2_1
XFILLER_106_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10210_ _10210_/A VGND VGND VPWR VPWR _11714_/A sky130_fd_sc_hd__inv_2
XFILLER_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11190_ _11190_/A VGND VGND VPWR VPWR _11190_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10141_ _10143_/A VGND VGND VPWR VPWR _10239_/B sky130_fd_sc_hd__buf_1
X_10072_ _10071_/A _10071_/B _09970_/A _10071_/X VGND VGND VPWR VPWR _10075_/A sky130_fd_sc_hd__a22o_1
X_13900_ _15414_/A _13955_/B VGND VGND VPWR VPWR _13900_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14880_ _14880_/A VGND VGND VPWR VPWR _15542_/A sky130_fd_sc_hd__buf_1
X_13831_ _14645_/A _13839_/B VGND VGND VPWR VPWR _13831_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13762_ _13762_/A _13762_/B VGND VGND VPWR VPWR _13762_/X sky130_fd_sc_hd__or2_1
XFILLER_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10974_ _10974_/A VGND VGND VPWR VPWR _10974_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15501_ _15449_/A _15449_/B _15449_/A _15449_/B VGND VGND VPWR VPWR _15501_/X sky130_fd_sc_hd__a2bb2o_1
X_12713_ _12699_/A _12699_/B _12699_/Y _12712_/X VGND VGND VPWR VPWR _12713_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13693_ _13738_/A _13691_/X _13692_/X VGND VGND VPWR VPWR _13693_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12644_ _12644_/A _12644_/B VGND VGND VPWR VPWR _12644_/Y sky130_fd_sc_hd__nand2_1
X_15432_ _15421_/Y _15431_/Y _15421_/Y _15431_/Y VGND VGND VPWR VPWR _15563_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12575_ _12624_/A _12624_/B VGND VGND VPWR VPWR _14213_/A sky130_fd_sc_hd__and2_1
X_15363_ _15363_/A _15349_/X VGND VGND VPWR VPWR _15363_/X sky130_fd_sc_hd__or2b_1
X_14314_ _14334_/A _14314_/B VGND VGND VPWR VPWR _15962_/A sky130_fd_sc_hd__or2_1
X_11526_ _11531_/A VGND VGND VPWR VPWR _11615_/A sky130_fd_sc_hd__inv_2
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15294_ _14833_/A _15237_/B _15237_/Y VGND VGND VPWR VPWR _15294_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14245_ _14361_/B VGND VGND VPWR VPWR _15781_/A sky130_fd_sc_hd__inv_2
X_11457_ _14113_/A _11386_/B _11386_/Y _12540_/A VGND VGND VPWR VPWR _12532_/A sky130_fd_sc_hd__a2bb2o_1
X_14176_ _14277_/A VGND VGND VPWR VPWR _15906_/A sky130_fd_sc_hd__buf_6
X_10408_ _10358_/X _10407_/X _10358_/X _10407_/X VGND VGND VPWR VPWR _10409_/B sky130_fd_sc_hd__a2bb2o_1
X_11388_ _08971_/X _11387_/X _08971_/X _11387_/X VGND VGND VPWR VPWR _11389_/B sky130_fd_sc_hd__a2bb2oi_2
X_13127_ _13984_/A _13127_/B VGND VGND VPWR VPWR _13127_/Y sky130_fd_sc_hd__nand2_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _09707_/A _09707_/B _09707_/Y VGND VGND VPWR VPWR _10339_/Y sky130_fd_sc_hd__a21oi_1
X_13058_ _13058_/A VGND VGND VPWR VPWR _13770_/A sky130_fd_sc_hd__inv_2
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12009_ _11984_/X _12008_/Y _11984_/X _12008_/Y VGND VGND VPWR VPWR _12070_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09220_ _09220_/A VGND VGND VPWR VPWR _09220_/Y sky130_fd_sc_hd__inv_2
X_09151_ _09518_/A _09148_/X _09148_/X _08524_/Y VGND VGND VPWR VPWR _09152_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09082_ _09763_/A VGND VGND VPWR VPWR _09436_/A sky130_fd_sc_hd__buf_1
XFILLER_116_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09984_ _09984_/A _09984_/B VGND VGND VPWR VPWR _09984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08935_ _08935_/A _08935_/B VGND VGND VPWR VPWR _08935_/X sky130_fd_sc_hd__or2_1
XFILLER_96_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08866_ _09486_/A _08776_/Y _08778_/Y _08865_/X VGND VGND VPWR VPWR _08866_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08797_ _08797_/A VGND VGND VPWR VPWR _08798_/A sky130_fd_sc_hd__inv_2
XFILLER_29_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10690_ _10678_/X _10689_/Y _10678_/X _10689_/Y VGND VGND VPWR VPWR _10812_/A sky130_fd_sc_hd__o2bb2a_1
X_09418_ _09418_/A _09418_/B VGND VGND VPWR VPWR _09418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09349_ _09527_/A _09743_/A VGND VGND VPWR VPWR _09350_/A sky130_fd_sc_hd__or2_1
X_12360_ _13204_/A _12360_/B VGND VGND VPWR VPWR _12360_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11311_ _11314_/A VGND VGND VPWR VPWR _11311_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12291_ _12255_/X _12290_/Y _12255_/X _12290_/Y VGND VGND VPWR VPWR _12360_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_107_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14030_ _13944_/X _14029_/Y _13944_/X _14029_/Y VGND VGND VPWR VPWR _14031_/B sky130_fd_sc_hd__a2bb2o_1
X_11242_ _11242_/A _11078_/X VGND VGND VPWR VPWR _11242_/X sky130_fd_sc_hd__or2b_1
XFILLER_134_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11173_ _11279_/A _11279_/B _11279_/A _11279_/B VGND VGND VPWR VPWR _11173_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10124_ _10124_/A _10124_/B VGND VGND VPWR VPWR _10125_/B sky130_fd_sc_hd__or2_1
X_15981_ _15982_/A _15982_/B VGND VGND VPWR VPWR _15981_/X sky130_fd_sc_hd__and2_1
XFILLER_79_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14932_ _15433_/A VGND VGND VPWR VPWR _15563_/A sky130_fd_sc_hd__buf_1
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10055_ _10055_/A _10055_/B VGND VGND VPWR VPWR _10055_/X sky130_fd_sc_hd__or2_1
X_14863_ _15552_/A _14928_/B VGND VGND VPWR VPWR _14863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13814_ _14618_/A _13849_/B VGND VGND VPWR VPWR _13814_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14794_ _14794_/A _14794_/B VGND VGND VPWR VPWR _14794_/X sky130_fd_sc_hd__and2_1
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13745_ _13687_/X _13744_/Y _13687_/X _13744_/Y VGND VGND VPWR VPWR _13758_/B sky130_fd_sc_hd__a2bb2o_1
X_10957_ _09990_/A _09990_/B _09990_/Y VGND VGND VPWR VPWR _10958_/A sky130_fd_sc_hd__o21ai_1
X_16464_ _16357_/A _16464_/D VGND VGND VPWR VPWR _16464_/Q sky130_fd_sc_hd__dfxtp_1
X_13676_ _13676_/A VGND VGND VPWR VPWR _14500_/A sky130_fd_sc_hd__inv_2
XFILLER_44_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12627_ _14207_/A _12625_/X _12626_/X VGND VGND VPWR VPWR _12627_/X sky130_fd_sc_hd__o21a_1
X_15415_ _15444_/A _15413_/X _15414_/X VGND VGND VPWR VPWR _15415_/X sky130_fd_sc_hd__o21a_1
X_10888_ _10888_/A VGND VGND VPWR VPWR _10888_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16395_ _16395_/A VGND VGND VPWR VPWR _16396_/B sky130_fd_sc_hd__inv_2
XFILLER_129_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12558_ _14914_/A _11449_/B _11449_/Y VGND VGND VPWR VPWR _12559_/A sky130_fd_sc_hd__o21ai_1
X_15346_ _15369_/A _15344_/X _15345_/X VGND VGND VPWR VPWR _15346_/X sky130_fd_sc_hd__o21a_1
X_12489_ _12486_/Y _12487_/Y _12488_/Y VGND VGND VPWR VPWR _12489_/Y sky130_fd_sc_hd__o21ai_1
X_15277_ _14581_/A _15255_/B _15255_/Y _15276_/X VGND VGND VPWR VPWR _15277_/X sky130_fd_sc_hd__a2bb2o_1
X_11509_ _11509_/A VGND VGND VPWR VPWR _13500_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14228_ _14906_/A _14083_/B _14083_/X VGND VGND VPWR VPWR _14228_/X sky130_fd_sc_hd__o21ba_1
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14159_ _13449_/A _14148_/B _14148_/Y VGND VGND VPWR VPWR _14159_/Y sky130_fd_sc_hd__a21oi_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08720_ _08856_/B VGND VGND VPWR VPWR _09540_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08651_ _08856_/B VGND VGND VPWR VPWR _08721_/B sky130_fd_sc_hd__inv_2
XFILLER_81_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08582_ _09454_/B VGND VGND VPWR VPWR _08714_/B sky130_fd_sc_hd__inv_2
XFILLER_50_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09203_ _11251_/B VGND VGND VPWR VPWR _11220_/B sky130_fd_sc_hd__buf_2
X_09134_ _09555_/B _09036_/B _09037_/B VGND VGND VPWR VPWR _09135_/A sky130_fd_sc_hd__a21bo_1
X_09065_ _09503_/B _09064_/A _09826_/B _09064_/Y VGND VGND VPWR VPWR _09069_/A sky130_fd_sc_hd__o22a_1
XFILLER_116_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09967_ _10081_/A VGND VGND VPWR VPWR _09967_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08918_ _09677_/A VGND VGND VPWR VPWR _08930_/A sky130_fd_sc_hd__inv_2
XFILLER_85_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09898_/A _09898_/B VGND VGND VPWR VPWR _09898_/X sky130_fd_sc_hd__and2_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08849_ _08935_/B VGND VGND VPWR VPWR _10103_/A sky130_fd_sc_hd__inv_2
XFILLER_72_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11860_ _10568_/A _11859_/A _10568_/Y _11923_/B VGND VGND VPWR VPWR _11862_/B sky130_fd_sc_hd__o22a_1
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11791_ _11791_/A VGND VGND VPWR VPWR _12830_/A sky130_fd_sc_hd__buf_1
X_10811_ _11992_/A VGND VGND VPWR VPWR _11928_/A sky130_fd_sc_hd__inv_2
XFILLER_26_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13530_ _12833_/A _12833_/B _10426_/B _12833_/Y VGND VGND VPWR VPWR _13530_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10742_ _09958_/A _09640_/B _09640_/Y VGND VGND VPWR VPWR _10744_/A sky130_fd_sc_hd__o21ai_1
X_15200_ _15134_/A _15134_/B _15134_/Y VGND VGND VPWR VPWR _15200_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10673_ _10675_/A VGND VGND VPWR VPWR _10673_/Y sky130_fd_sc_hd__inv_2
X_13461_ _11612_/Y _12678_/X _11694_/X VGND VGND VPWR VPWR _13461_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16180_ _16107_/X _16179_/X _16107_/X _16179_/X VGND VGND VPWR VPWR _16181_/B sky130_fd_sc_hd__a2bb2oi_1
X_13392_ _14113_/A _13437_/B VGND VGND VPWR VPWR _13392_/Y sky130_fd_sc_hd__nor2_1
X_12412_ _12412_/A _12412_/B VGND VGND VPWR VPWR _12412_/Y sky130_fd_sc_hd__nand2_1
X_12343_ _12346_/A _12346_/B VGND VGND VPWR VPWR _12343_/Y sky130_fd_sc_hd__nor2_1
X_15131_ _15131_/A _15131_/B VGND VGND VPWR VPWR _15131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15062_ _15041_/X _15061_/X _15041_/X _15061_/X VGND VGND VPWR VPWR _15063_/B sky130_fd_sc_hd__a2bb2o_1
X_12274_ _12275_/A _12275_/B VGND VGND VPWR VPWR _12274_/X sky130_fd_sc_hd__and2_1
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11225_ _14031_/A _11225_/B VGND VGND VPWR VPWR _11225_/Y sky130_fd_sc_hd__nand2_1
X_14013_ _13954_/X _14012_/Y _13954_/X _14012_/Y VGND VGND VPWR VPWR _14059_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11156_ _11155_/A _11155_/B _11155_/Y _10984_/X VGND VGND VPWR VPWR _12268_/A sky130_fd_sc_hd__o211a_1
X_15964_ _15964_/A _15964_/B VGND VGND VPWR VPWR _15999_/B sky130_fd_sc_hd__or2_1
X_11087_ _11217_/A _11085_/X _11086_/X VGND VGND VPWR VPWR _11087_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10107_ _10177_/A _10177_/B _10106_/Y VGND VGND VPWR VPWR _10109_/A sky130_fd_sc_hd__o21ai_1
X_14915_ _14889_/Y _14913_/X _14914_/Y VGND VGND VPWR VPWR _14915_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10038_ _10038_/A _10038_/B VGND VGND VPWR VPWR _10038_/Y sky130_fd_sc_hd__nor2_1
X_15895_ _15871_/Y _15893_/X _15894_/Y VGND VGND VPWR VPWR _15895_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14846_ _14837_/X _14845_/Y _14837_/X _14845_/Y VGND VGND VPWR VPWR _14848_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14777_ _14739_/X _14776_/X _14739_/X _14776_/X VGND VGND VPWR VPWR _14778_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13728_ _13770_/A _13770_/B VGND VGND VPWR VPWR _13806_/A sky130_fd_sc_hd__and2_1
X_11989_ _11987_/A _11987_/B _11987_/X _11988_/Y VGND VGND VPWR VPWR _12077_/B sky130_fd_sc_hd__a22o_1
XFILLER_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16447_ _16447_/A _16447_/B VGND VGND VPWR VPWR _16447_/X sky130_fd_sc_hd__or2_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13659_ _13635_/A _13658_/Y _13635_/A _13658_/Y VGND VGND VPWR VPWR _13698_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16378_ _16318_/A _16318_/B _16318_/Y VGND VGND VPWR VPWR _16378_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15329_ _15329_/A _15329_/B VGND VGND VPWR VPWR _15329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09821_ _09821_/A _09821_/B VGND VGND VPWR VPWR _09882_/B sky130_fd_sc_hd__or2_1
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09752_ _10087_/A VGND VGND VPWR VPWR _09997_/B sky130_fd_sc_hd__buf_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _08703_/A VGND VGND VPWR VPWR _09937_/A sky130_fd_sc_hd__inv_2
XFILLER_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09683_ _09683_/A _09683_/B VGND VGND VPWR VPWR _09686_/A sky130_fd_sc_hd__or2_1
XFILLER_27_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08634_ _08634_/A VGND VGND VPWR VPWR _09462_/B sky130_fd_sc_hd__inv_2
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08565_ _10012_/A _08565_/B VGND VGND VPWR VPWR _09858_/A sky130_fd_sc_hd__or2_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08496_ _08239_/Y _08699_/A _08237_/A _08235_/B VGND VGND VPWR VPWR _08496_/X sky130_fd_sc_hd__o22a_2
XFILLER_23_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09117_ _09117_/A VGND VGND VPWR VPWR _09117_/Y sky130_fd_sc_hd__inv_2
X_09048_ _08714_/Y _09047_/Y _08730_/X VGND VGND VPWR VPWR _09048_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11010_ _13583_/A VGND VGND VPWR VPWR _12853_/A sky130_fd_sc_hd__buf_1
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12961_ _14757_/A _12946_/B _12946_/Y VGND VGND VPWR VPWR _12961_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15680_ _15607_/Y _15678_/X _15679_/Y VGND VGND VPWR VPWR _15680_/X sky130_fd_sc_hd__o21a_1
X_14700_ _14654_/X _14699_/Y _14654_/X _14699_/Y VGND VGND VPWR VPWR _14732_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12892_ _14468_/A _12936_/B VGND VGND VPWR VPWR _12892_/Y sky130_fd_sc_hd__nor2_1
X_11912_ _13632_/A _11912_/B VGND VGND VPWR VPWR _11912_/Y sky130_fd_sc_hd__nor2_1
X_14631_ _14577_/A _14577_/B _14577_/Y VGND VGND VPWR VPWR _14631_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11843_ _11827_/Y _11841_/X _11842_/Y VGND VGND VPWR VPWR _11843_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16301_ _16256_/X _16300_/Y _16256_/X _16300_/Y VGND VGND VPWR VPWR _16324_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14575_/A _14575_/B VGND VGND VPWR VPWR _14562_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11774_ _11774_/A VGND VGND VPWR VPWR _12768_/A sky130_fd_sc_hd__buf_1
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _14462_/A _14462_/B _14462_/Y VGND VGND VPWR VPWR _14493_/Y sky130_fd_sc_hd__o21ai_1
X_13513_ _13515_/A VGND VGND VPWR VPWR _15038_/A sky130_fd_sc_hd__buf_1
XFILLER_9_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10725_ _09975_/A _09650_/B _09650_/Y VGND VGND VPWR VPWR _10727_/A sky130_fd_sc_hd__o21ai_1
X_16232_ _16084_/A _16084_/B _16084_/Y VGND VGND VPWR VPWR _16234_/A sky130_fd_sc_hd__o21ai_1
X_13444_ _13383_/Y _13442_/X _13443_/Y VGND VGND VPWR VPWR _13444_/X sky130_fd_sc_hd__o21a_1
X_10656_ _10656_/A VGND VGND VPWR VPWR _10656_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16163_ _16070_/X _16163_/B VGND VGND VPWR VPWR _16163_/X sky130_fd_sc_hd__and2b_1
XFILLER_70_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13375_ _13313_/A _13313_/B _13313_/A _13313_/B VGND VGND VPWR VPWR _13375_/X sky130_fd_sc_hd__a2bb2o_1
X_15114_ _15057_/A _15057_/B _15057_/Y VGND VGND VPWR VPWR _15114_/Y sky130_fd_sc_hd__o21ai_1
X_10587_ _09970_/Y _10586_/A _09970_/A _10586_/Y _10943_/A VGND VGND VPWR VPWR _11907_/A
+ sky130_fd_sc_hd__a221o_2
X_16094_ _16094_/A _16094_/B VGND VGND VPWR VPWR _16094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12326_ _12239_/X _12325_/Y _12239_/X _12325_/Y VGND VGND VPWR VPWR _12601_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12257_ _12257_/A VGND VGND VPWR VPWR _12257_/Y sky130_fd_sc_hd__inv_2
X_15045_ _15058_/A _15043_/X _15044_/X VGND VGND VPWR VPWR _15045_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11208_ _13331_/A VGND VGND VPWR VPWR _12217_/A sky130_fd_sc_hd__inv_2
X_12188_ _12168_/X _12187_/X _12168_/X _12187_/X VGND VGND VPWR VPWR _12259_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11139_ _11136_/Y _12689_/A _10965_/X _11138_/Y VGND VGND VPWR VPWR _11139_/X sky130_fd_sc_hd__o22a_1
X_15947_ _15947_/A _15947_/B VGND VGND VPWR VPWR _15947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15878_ _15878_/A VGND VGND VPWR VPWR _15888_/A sky130_fd_sc_hd__inv_2
XFILLER_76_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14829_ _14741_/X _14772_/A _14771_/X VGND VGND VPWR VPWR _14829_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08350_ _08348_/Y _08349_/A _08348_/A _08349_/Y _08303_/A VGND VGND VPWR VPWR _09221_/B
+ sky130_fd_sc_hd__o221a_1
X_08281_ _08358_/A input18/X VGND VGND VPWR VPWR _08282_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ _09856_/B VGND VGND VPWR VPWR _09804_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09735_ _08558_/A _09737_/B _08558_/A _09737_/B VGND VGND VPWR VPWR _09736_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09666_ _09997_/A _09666_/B VGND VGND VPWR VPWR _09666_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08617_ _08716_/A VGND VGND VPWR VPWR _09456_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09597_ _09987_/A _09658_/B VGND VGND VPWR VPWR _09597_/Y sky130_fd_sc_hd__nor2_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08690_/A _10118_/B VGND VGND VPWR VPWR _08881_/A sky130_fd_sc_hd__nor2_1
X_08479_ input27/X input11/X VGND VGND VPWR VPWR _08479_/Y sky130_fd_sc_hd__nor2_1
X_10510_ _11838_/A VGND VGND VPWR VPWR _15143_/A sky130_fd_sc_hd__buf_1
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11490_ _09665_/X _11489_/X _09665_/X _11489_/X VGND VGND VPWR VPWR _11491_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_109_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10441_ _13521_/A _10441_/B VGND VGND VPWR VPWR _10441_/X sky130_fd_sc_hd__and2_1
XFILLER_7_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13160_ _15252_/A _13113_/B _13113_/Y VGND VGND VPWR VPWR _13160_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10372_ _09117_/A _10371_/X _09117_/A _10371_/X VGND VGND VPWR VPWR _11220_/A sky130_fd_sc_hd__a2bb2o_2
X_12111_ _12064_/X _12110_/Y _12064_/X _12110_/Y VGND VGND VPWR VPWR _12153_/B sky130_fd_sc_hd__a2bb2o_1
X_13091_ _13013_/X _13090_/X _13013_/X _13090_/X VGND VGND VPWR VPWR _13105_/B sky130_fd_sc_hd__a2bb2o_1
X_12042_ _13184_/A _12051_/B VGND VGND VPWR VPWR _12042_/Y sky130_fd_sc_hd__nor2_1
X_15801_ _15797_/Y _16217_/A _15800_/Y VGND VGND VPWR VPWR _15805_/B sky130_fd_sc_hd__o21ai_1
X_13993_ _15422_/A _13994_/B VGND VGND VPWR VPWR _13993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15732_ _15544_/A _14920_/B _14920_/Y VGND VGND VPWR VPWR _15732_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12944_ _12944_/A _12944_/B VGND VGND VPWR VPWR _12944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15663_ _15947_/A _15662_/B _14374_/A _14374_/Y _15662_/Y VGND VGND VPWR VPWR _15665_/B
+ sky130_fd_sc_hd__o32a_1
X_12875_ _12856_/X _12874_/Y _12856_/X _12874_/Y VGND VGND VPWR VPWR _12944_/B sky130_fd_sc_hd__a2bb2o_1
X_15594_ _15543_/X _15593_/X _15543_/X _15593_/X VGND VGND VPWR VPWR _15595_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14614_/A VGND VGND VPWR VPWR _15343_/A sky130_fd_sc_hd__buf_1
X_11826_ _11798_/X _11825_/X _11798_/X _11825_/X VGND VGND VPWR VPWR _11842_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14518_/X _14544_/X _14518_/X _14544_/X VGND VGND VPWR VPWR _14583_/B sky130_fd_sc_hd__a2bb2o_1
X_11757_ _11774_/A _11744_/B _11744_/X _11756_/Y VGND VGND VPWR VPWR _11801_/B sky130_fd_sc_hd__a22o_1
XFILLER_81_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10708_ _11942_/A _10708_/B VGND VGND VPWR VPWR _10708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16215_ _16213_/A _16214_/A _16213_/Y _16214_/Y _16205_/A VGND VGND VPWR VPWR _16253_/A
+ sky130_fd_sc_hd__a221o_1
X_11688_ _11688_/A VGND VGND VPWR VPWR _11688_/Y sky130_fd_sc_hd__inv_2
X_14476_ _14476_/A _14476_/B VGND VGND VPWR VPWR _14476_/Y sky130_fd_sc_hd__nor2_1
X_13427_ _14105_/A _13430_/B VGND VGND VPWR VPWR _13427_/Y sky130_fd_sc_hd__nor2_1
X_10639_ _12992_/A _10639_/B VGND VGND VPWR VPWR _10639_/Y sky130_fd_sc_hd__nand2_1
X_16146_ _16119_/A _16119_/B _16119_/Y VGND VGND VPWR VPWR _16148_/A sky130_fd_sc_hd__o21ai_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13358_ _13340_/A _13340_/B _13340_/X _13357_/X VGND VGND VPWR VPWR _13358_/X sky130_fd_sc_hd__o22a_1
X_16077_ _16038_/A _16038_/B _16038_/Y VGND VGND VPWR VPWR _16077_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_115_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12309_ _14017_/A _12211_/B _12211_/Y VGND VGND VPWR VPWR _12309_/Y sky130_fd_sc_hd__o21ai_1
X_13289_ _13245_/Y _13287_/Y _13288_/Y VGND VGND VPWR VPWR _13290_/A sky130_fd_sc_hd__o21ai_1
X_15028_ _15028_/A _15028_/B VGND VGND VPWR VPWR _15028_/X sky130_fd_sc_hd__or2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 wbs_adr_i[10] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_2
X_09520_ _09340_/A _08706_/B _09520_/S VGND VGND VPWR VPWR _09520_/X sky130_fd_sc_hd__mux2_1
X_09451_ _09486_/A _09529_/A VGND VGND VPWR VPWR _09451_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09382_ _09432_/B _09382_/B VGND VGND VPWR VPWR _09382_/X sky130_fd_sc_hd__or2_1
X_08402_ _08670_/A VGND VGND VPWR VPWR _08402_/X sky130_fd_sc_hd__clkbuf_2
X_08333_ _08333_/A VGND VGND VPWR VPWR _08333_/Y sky130_fd_sc_hd__inv_2
X_08264_ input13/X VGND VGND VPWR VPWR _08346_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_32_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09718_ _09963_/A _10597_/A _09717_/X VGND VGND VPWR VPWR _09720_/B sky130_fd_sc_hd__o21ai_1
X_10990_ _13506_/A _11130_/B _13506_/A _11130_/B VGND VGND VPWR VPWR _10990_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09649_ _09648_/A _09648_/B _09546_/A _09546_/Y _09648_/Y VGND VGND VPWR VPWR _10726_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_82_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12660_ _10369_/Y _12659_/Y _10307_/Y VGND VGND VPWR VPWR _12661_/A sky130_fd_sc_hd__o21ai_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11611_ _10122_/Y _11610_/A _10237_/B _11610_/Y _11529_/A VGND VGND VPWR VPWR _12426_/B
+ sky130_fd_sc_hd__a221o_1
X_14330_ _15869_/A _14262_/B _14262_/Y VGND VGND VPWR VPWR _14330_/Y sky130_fd_sc_hd__o21ai_1
X_12591_ _12591_/A _12331_/X VGND VGND VPWR VPWR _12592_/A sky130_fd_sc_hd__or2b_1
X_11542_ _11511_/X _11541_/X _11511_/X _11541_/X VGND VGND VPWR VPWR _11634_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14261_ _14261_/A VGND VGND VPWR VPWR _14261_/Y sky130_fd_sc_hd__inv_2
X_11473_ _14005_/A VGND VGND VPWR VPWR _14065_/A sky130_fd_sc_hd__buf_1
XFILLER_11_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16000_ _15963_/X _15999_/Y _15963_/X _15999_/Y VGND VGND VPWR VPWR _16046_/B sky130_fd_sc_hd__a2bb2o_1
X_14192_ _13437_/A _14114_/A _14078_/Y VGND VGND VPWR VPWR _14192_/Y sky130_fd_sc_hd__a21oi_1
X_13212_ _14841_/A VGND VGND VPWR VPWR _14858_/A sky130_fd_sc_hd__buf_1
X_10424_ _10424_/A _10424_/B VGND VGND VPWR VPWR _10425_/A sky130_fd_sc_hd__or2_1
X_13143_ _13124_/X _13142_/Y _13124_/X _13142_/Y VGND VGND VPWR VPWR _13206_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_97_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10355_ _12832_/A _10355_/B VGND VGND VPWR VPWR _10356_/A sky130_fd_sc_hd__nand2_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13074_ _13764_/A VGND VGND VPWR VPWR _15255_/A sky130_fd_sc_hd__buf_1
X_10286_ _13478_/A _10286_/B VGND VGND VPWR VPWR _10289_/A sky130_fd_sc_hd__and2_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12025_ _12059_/A VGND VGND VPWR VPWR _13192_/A sky130_fd_sc_hd__buf_1
XFILLER_78_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13976_ _13973_/X _13997_/A _13973_/X _13997_/A VGND VGND VPWR VPWR _13978_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15715_ _15728_/A _15715_/B VGND VGND VPWR VPWR _16121_/A sky130_fd_sc_hd__or2_1
XFILLER_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12927_ _12912_/Y _12924_/Y _12926_/Y VGND VGND VPWR VPWR _12927_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15646_ _15669_/A _15669_/B VGND VGND VPWR VPWR _15646_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12858_ _12799_/Y _12856_/X _12857_/Y VGND VGND VPWR VPWR _12858_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11809_ _10374_/A _11764_/A _10452_/B _11808_/Y VGND VGND VPWR VPWR _11810_/A sky130_fd_sc_hd__o22a_1
XFILLER_21_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15577_ _14401_/X _15576_/Y _14401_/X _15576_/Y VGND VGND VPWR VPWR _15696_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12789_ _12789_/A _12789_/B VGND VGND VPWR VPWR _12789_/Y sky130_fd_sc_hd__nor2_1
X_14528_ _14528_/A _14528_/B VGND VGND VPWR VPWR _14528_/Y sky130_fd_sc_hd__nor2_1
X_14459_ _14456_/Y _14457_/Y _14458_/Y VGND VGND VPWR VPWR _14459_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16129_ _15987_/X _16128_/X _15987_/X _16128_/X VGND VGND VPWR VPWR _16243_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_130_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08951_ _08680_/X _08950_/Y _08680_/X _08950_/Y VGND VGND VPWR VPWR _08951_/Y sky130_fd_sc_hd__a2bb2oi_2
X_08882_ _08689_/X _08881_/Y _08689_/X _08881_/Y VGND VGND VPWR VPWR _08980_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09503_ _09503_/A _09503_/B VGND VGND VPWR VPWR _09503_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09434_ _09247_/A _09433_/Y _09426_/Y VGND VGND VPWR VPWR _09436_/B sky130_fd_sc_hd__o21ai_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09365_ _09476_/B _09862_/A _09348_/A VGND VGND VPWR VPWR _09365_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09296_ _09296_/A VGND VGND VPWR VPWR _09296_/Y sky130_fd_sc_hd__inv_2
X_08316_ _08316_/A input20/X VGND VGND VPWR VPWR _08317_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08247_ input20/X VGND VGND VPWR VPWR _08248_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10140_ _10119_/A _10119_/B _10120_/A VGND VGND VPWR VPWR _10143_/A sky130_fd_sc_hd__a21bo_1
XFILLER_102_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10071_ _10071_/A _10071_/B VGND VGND VPWR VPWR _10071_/X sky130_fd_sc_hd__or2_1
XFILLER_48_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13830_ _13755_/X _13829_/Y _13755_/X _13829_/Y VGND VGND VPWR VPWR _13839_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13761_ _13821_/A _13759_/X _13760_/X VGND VGND VPWR VPWR _13761_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10973_ _10241_/B _10151_/B _10151_/Y VGND VGND VPWR VPWR _10974_/A sky130_fd_sc_hd__a21oi_1
X_15500_ _15546_/A _15546_/B VGND VGND VPWR VPWR _15500_/X sky130_fd_sc_hd__and2_1
XFILLER_90_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12712_ _12701_/A _12701_/B _12701_/Y _12711_/X VGND VGND VPWR VPWR _12712_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15431_ _15422_/A _15422_/B _15422_/Y VGND VGND VPWR VPWR _15431_/Y sky130_fd_sc_hd__o21ai_1
X_13692_ _13692_/A _13692_/B VGND VGND VPWR VPWR _13692_/X sky130_fd_sc_hd__or2_1
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12643_ _11674_/X _12643_/B VGND VGND VPWR VPWR _12644_/B sky130_fd_sc_hd__and2b_1
XFILLER_62_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12574_ _12571_/Y _12573_/Y _12571_/A _12573_/A _12503_/A VGND VGND VPWR VPWR _12624_/B
+ sky130_fd_sc_hd__o221a_1
X_15362_ _15418_/A _15418_/B VGND VGND VPWR VPWR _15362_/X sky130_fd_sc_hd__and2_1
XFILLER_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14313_ _13438_/X _14312_/X _13438_/X _14312_/X VGND VGND VPWR VPWR _14314_/B sky130_fd_sc_hd__a2bb2oi_1
X_15293_ _15353_/A _15353_/B VGND VGND VPWR VPWR _15293_/X sky130_fd_sc_hd__and2_1
X_11525_ _11607_/A _11525_/B VGND VGND VPWR VPWR _11531_/A sky130_fd_sc_hd__or2_1
XFILLER_7_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14244_ _14244_/A _14361_/B VGND VGND VPWR VPWR _14247_/A sky130_fd_sc_hd__or2_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11456_ _11451_/Y _12546_/A _11455_/Y VGND VGND VPWR VPWR _12540_/A sky130_fd_sc_hd__o21ai_2
XFILLER_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14175_ _14281_/A _14175_/B VGND VGND VPWR VPWR _14277_/A sky130_fd_sc_hd__or2_1
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10407_ _13527_/A _10328_/B _10324_/A _10328_/B VGND VGND VPWR VPWR _10407_/X sky130_fd_sc_hd__a2bb2o_1
X_11387_ _08907_/X _11387_/B VGND VGND VPWR VPWR _11387_/X sky130_fd_sc_hd__and2b_1
X_13126_ _13042_/Y _13124_/X _13125_/Y VGND VGND VPWR VPWR _13126_/X sky130_fd_sc_hd__o21a_1
X_10338_ _13529_/A _10338_/B VGND VGND VPWR VPWR _10338_/X sky130_fd_sc_hd__and2_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13057_ _15243_/A _13119_/B VGND VGND VPWR VPWR _13057_/Y sky130_fd_sc_hd__nor2_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12008_ _12007_/A _12073_/B _12007_/Y VGND VGND VPWR VPWR _12008_/Y sky130_fd_sc_hd__o21ai_1
X_10269_ _10234_/Y _10235_/X _10175_/Y _10236_/Y _10471_/A VGND VGND VPWR VPWR _11745_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13959_ _15418_/A _13959_/B VGND VGND VPWR VPWR _13959_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15629_ _14382_/X _15628_/Y _14382_/X _15628_/Y VGND VGND VPWR VPWR _15673_/B sky130_fd_sc_hd__a2bb2o_1
X_09150_ _08512_/X _09146_/X _09150_/S VGND VGND VPWR VPWR _09561_/B sky130_fd_sc_hd__mux2_1
X_09081_ _10012_/B _09077_/B _09078_/B VGND VGND VPWR VPWR _09763_/A sky130_fd_sc_hd__a21bo_1
XFILLER_131_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09983_ _09983_/A _09984_/B VGND VGND VPWR VPWR _09983_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08934_ _08934_/A VGND VGND VPWR VPWR _08935_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08865_ _09488_/A _08784_/Y _08786_/Y _08864_/X VGND VGND VPWR VPWR _08865_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08796_ _09209_/A _09453_/B _08713_/X VGND VGND VPWR VPWR _08797_/A sky130_fd_sc_hd__o21ai_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09417_ _09418_/A _09418_/B VGND VGND VPWR VPWR _09417_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09348_ _09348_/A VGND VGND VPWR VPWR _09348_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09279_ _08623_/A _09802_/A _09224_/A VGND VGND VPWR VPWR _09279_/X sky130_fd_sc_hd__o21a_1
X_11310_ _11309_/A _11309_/B _11309_/Y _10959_/X VGND VGND VPWR VPWR _11509_/A sky130_fd_sc_hd__o211a_1
XFILLER_119_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12290_ _12289_/A _12362_/B _12289_/Y VGND VGND VPWR VPWR _12290_/Y sky130_fd_sc_hd__o21ai_1
X_11241_ _12232_/A VGND VGND VPWR VPWR _13348_/A sky130_fd_sc_hd__buf_1
XFILLER_4_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11172_ _11110_/X _11171_/Y _11110_/X _11171_/Y VGND VGND VPWR VPWR _11279_/B sky130_fd_sc_hd__o2bb2a_1
X_10123_ _10123_/A _10123_/B VGND VGND VPWR VPWR _10124_/B sky130_fd_sc_hd__or2_1
X_15980_ _15977_/Y _15979_/X _15977_/Y _15979_/X VGND VGND VPWR VPWR _15982_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14931_ _14930_/A _14930_/B _14827_/X _14930_/X VGND VGND VPWR VPWR _14931_/X sky130_fd_sc_hd__o22a_1
X_10054_ _08930_/A _09505_/Y _08916_/A _09505_/A VGND VGND VPWR VPWR _10055_/B sky130_fd_sc_hd__o22a_1
X_14862_ _14827_/X _14861_/X _14827_/X _14861_/X VGND VGND VPWR VPWR _14928_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13813_ _13765_/X _13812_/X _13765_/X _13812_/X VGND VGND VPWR VPWR _13849_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14793_ _14731_/X _14792_/X _14731_/X _14792_/X VGND VGND VPWR VPWR _14794_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13744_ _14496_/A _13688_/B _13688_/Y VGND VGND VPWR VPWR _13744_/Y sky130_fd_sc_hd__o21ai_1
X_10956_ _13509_/A _10955_/B _10955_/X _10805_/X VGND VGND VPWR VPWR _10956_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16463_ _16357_/A _16463_/D VGND VGND VPWR VPWR _16463_/Q sky130_fd_sc_hd__dfxtp_1
X_13675_ _14496_/A _13688_/B VGND VGND VPWR VPWR _13675_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10887_ _09409_/A _09409_/B _09409_/Y VGND VGND VPWR VPWR _10888_/A sky130_fd_sc_hd__a21oi_1
XFILLER_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16394_ _16407_/C _16407_/A VGND VGND VPWR VPWR _16394_/Y sky130_fd_sc_hd__nand2_1
X_12626_ _12626_/A _12626_/B VGND VGND VPWR VPWR _12626_/X sky130_fd_sc_hd__or2_1
X_15414_ _15414_/A _15414_/B VGND VGND VPWR VPWR _15414_/X sky130_fd_sc_hd__or2_1
X_15345_ _15345_/A _15345_/B VGND VGND VPWR VPWR _15345_/X sky130_fd_sc_hd__or2_1
XFILLER_12_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12557_ _15534_/A VGND VGND VPWR VPWR _14914_/A sky130_fd_sc_hd__buf_1
XFILLER_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12488_ _13132_/A _12488_/B VGND VGND VPWR VPWR _12488_/Y sky130_fd_sc_hd__nand2_1
X_15276_ _14579_/A _15258_/B _15258_/Y _15275_/X VGND VGND VPWR VPWR _15276_/X sky130_fd_sc_hd__a2bb2o_1
X_11508_ _12442_/A VGND VGND VPWR VPWR _13871_/A sky130_fd_sc_hd__buf_1
X_14227_ _15878_/A _14253_/B VGND VGND VPWR VPWR _14227_/Y sky130_fd_sc_hd__nor2_1
X_11439_ _13395_/A _11443_/B VGND VGND VPWR VPWR _11439_/Y sky130_fd_sc_hd__nor2_1
X_14158_ _14206_/A VGND VGND VPWR VPWR _14281_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13109_ _15258_/A _13109_/B VGND VGND VPWR VPWR _13109_/Y sky130_fd_sc_hd__nand2_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14089_ _14049_/X _14088_/X _14049_/X _14088_/X VGND VGND VPWR VPWR _14089_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08650_ _08650_/A _08650_/B VGND VGND VPWR VPWR _08856_/B sky130_fd_sc_hd__or2_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08581_ _08580_/X _08428_/X _08580_/X _08428_/X VGND VGND VPWR VPWR _08584_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09202_ _11413_/B VGND VGND VPWR VPWR _11251_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09133_ _09426_/A _09136_/B VGND VGND VPWR VPWR _09133_/Y sky130_fd_sc_hd__nor2_1
X_09064_ _09064_/A VGND VGND VPWR VPWR _09064_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09966_ _10083_/A VGND VGND VPWR VPWR _09966_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09854_/B _09897_/B VGND VGND VPWR VPWR _09898_/B sky130_fd_sc_hd__nand2b_1
X_08917_ _08917_/A VGND VGND VPWR VPWR _08922_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _09503_/B _08722_/X _08847_/A _08722_/X VGND VGND VPWR VPWR _08935_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08779_ _09452_/A VGND VGND VPWR VPWR _09488_/A sky130_fd_sc_hd__buf_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11790_ _11790_/A _11790_/B VGND VGND VPWR VPWR _11790_/Y sky130_fd_sc_hd__nor2_1
X_10810_ _10812_/A VGND VGND VPWR VPWR _10810_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10741_ _11970_/A _10741_/B VGND VGND VPWR VPWR _10741_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13460_ _15425_/A _12864_/B _12864_/Y _12950_/X VGND VGND VPWR VPWR _13460_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12411_ _13447_/A _12410_/B _12410_/Y VGND VGND VPWR VPWR _12412_/B sky130_fd_sc_hd__o21a_1
X_10672_ _11919_/A VGND VGND VPWR VPWR _13512_/A sky130_fd_sc_hd__buf_1
XFILLER_43_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13391_ _13361_/X _13390_/X _13361_/X _13390_/X VGND VGND VPWR VPWR _13437_/B sky130_fd_sc_hd__a2bb2o_1
X_12342_ _12338_/Y _12571_/A _12341_/Y VGND VGND VPWR VPWR _12346_/B sky130_fd_sc_hd__o21ai_1
X_15130_ _15092_/X _15129_/Y _15092_/X _15129_/Y VGND VGND VPWR VPWR _15131_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15061_ _15061_/A _15042_/X VGND VGND VPWR VPWR _15061_/X sky130_fd_sc_hd__or2b_1
X_12273_ _11328_/A _12272_/A _11328_/Y _12272_/Y VGND VGND VPWR VPWR _12275_/B sky130_fd_sc_hd__o22a_1
XFILLER_5_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14012_ _15414_/A _13955_/B _13955_/Y VGND VGND VPWR VPWR _14012_/Y sky130_fd_sc_hd__o21ai_1
X_11224_ _11083_/X _11223_/X _11083_/X _11223_/X VGND VGND VPWR VPWR _11225_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11155_ _11155_/A _11155_/B VGND VGND VPWR VPWR _11155_/Y sky130_fd_sc_hd__nand2_1
X_15963_ _15924_/X _15961_/X _16002_/B VGND VGND VPWR VPWR _15963_/X sky130_fd_sc_hd__o21a_1
X_11086_ _13913_/A _11086_/B VGND VGND VPWR VPWR _11086_/X sky130_fd_sc_hd__or2_1
X_10106_ _10177_/A _10177_/B VGND VGND VPWR VPWR _10106_/Y sky130_fd_sc_hd__nand2_1
X_14914_ _14914_/A _14914_/B VGND VGND VPWR VPWR _14914_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10037_ _10087_/A _10087_/B VGND VGND VPWR VPWR _10037_/X sky130_fd_sc_hd__and2_1
XFILLER_124_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15894_ _15894_/A _15894_/B VGND VGND VPWR VPWR _15894_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14845_ _14944_/A _14944_/B _14844_/Y VGND VGND VPWR VPWR _14845_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14776_ _14776_/A _14740_/X VGND VGND VPWR VPWR _14776_/X sky130_fd_sc_hd__or2b_1
X_11988_ _11988_/A VGND VGND VPWR VPWR _11988_/Y sky130_fd_sc_hd__inv_2
X_13727_ _13699_/X _13726_/X _13699_/X _13726_/X VGND VGND VPWR VPWR _13770_/B sky130_fd_sc_hd__a2bb2o_1
X_10939_ _10939_/A VGND VGND VPWR VPWR _10939_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16446_ _16471_/Q VGND VGND VPWR VPWR _16446_/Y sky130_fd_sc_hd__inv_2
X_13658_ _15125_/A _13637_/B _13637_/Y VGND VGND VPWR VPWR _13658_/Y sky130_fd_sc_hd__o21ai_1
X_16377_ _08230_/A _16460_/Q _08233_/A _16397_/A _16343_/A VGND VGND VPWR VPWR _16460_/D
+ sky130_fd_sc_hd__o221a_2
X_12609_ _14243_/A _12608_/B _12608_/Y _11708_/A VGND VGND VPWR VPWR _14234_/A sky130_fd_sc_hd__o211a_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13589_ _13636_/A _13637_/B VGND VGND VPWR VPWR _13589_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15328_ _11066_/B _15327_/X _11066_/B _15327_/X VGND VGND VPWR VPWR _15329_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15259_ _15205_/A _15205_/B _15205_/Y VGND VGND VPWR VPWR _15259_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09820_ _09820_/A _09820_/B VGND VGND VPWR VPWR _09821_/B sky130_fd_sc_hd__or2_1
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09751_ _09745_/A _09745_/B _09791_/A VGND VGND VPWR VPWR _10087_/A sky130_fd_sc_hd__a21bo_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ _08703_/A _09146_/A VGND VGND VPWR VPWR _09340_/A sky130_fd_sc_hd__nor2_1
XFILLER_94_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09682_ _08657_/A _09684_/B _08657_/A _09684_/B VGND VGND VPWR VPWR _09683_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08633_ _08632_/X _08408_/Y _08632_/X _08408_/Y VGND VGND VPWR VPWR _08635_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _09453_/B VGND VGND VPWR VPWR _09555_/A sky130_fd_sc_hd__buf_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08495_ _08242_/A _08306_/B _08469_/Y _08501_/A VGND VGND VPWR VPWR _08699_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09116_ _09547_/B _09032_/B _09033_/B VGND VGND VPWR VPWR _09117_/A sky130_fd_sc_hd__a21bo_1
XFILLER_108_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09047_ _09047_/A VGND VGND VPWR VPWR _09047_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09949_ _09949_/A VGND VGND VPWR VPWR _11773_/A sky130_fd_sc_hd__buf_1
XFILLER_49_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12960_ _13792_/A VGND VGND VPWR VPWR _14749_/A sky130_fd_sc_hd__inv_2
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11911_ _11873_/Y _11909_/Y _11910_/Y VGND VGND VPWR VPWR _11981_/A sky130_fd_sc_hd__o21ai_1
X_12891_ _12848_/X _12890_/Y _12848_/X _12890_/Y VGND VGND VPWR VPWR _12936_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14630_/A VGND VGND VPWR VPWR _15335_/A sky130_fd_sc_hd__buf_1
X_11842_ _11842_/A _11842_/B VGND VGND VPWR VPWR _11842_/Y sky130_fd_sc_hd__nand2_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14510_/X _14560_/X _14510_/X _14560_/X VGND VGND VPWR VPWR _14575_/B sky130_fd_sc_hd__a2bb2o_1
X_16300_ _16324_/A _16258_/B _16258_/Y VGND VGND VPWR VPWR _16300_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11773_/A _11773_/B VGND VGND VPWR VPWR _11773_/X sky130_fd_sc_hd__and2_1
X_13512_ _13512_/A _13512_/B VGND VGND VPWR VPWR _13512_/Y sky130_fd_sc_hd__nand2_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14492_/A VGND VGND VPWR VPWR _15205_/A sky130_fd_sc_hd__buf_1
X_10724_ _13073_/A _10724_/B VGND VGND VPWR VPWR _10724_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16231_ _16251_/A _16318_/A VGND VGND VPWR VPWR _16231_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13443_ _13443_/A _13443_/B VGND VGND VPWR VPWR _13443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10655_ _10654_/Y _10534_/X _10581_/Y VGND VGND VPWR VPWR _10655_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16162_ _16268_/A _16334_/A VGND VGND VPWR VPWR _16162_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13374_ _13449_/A _13449_/B VGND VGND VPWR VPWR _13374_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12325_ _12232_/A _12232_/B _12232_/Y VGND VGND VPWR VPWR _12325_/Y sky130_fd_sc_hd__o21ai_1
X_15113_ _15113_/A _15113_/B VGND VGND VPWR VPWR _15113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10586_ _10586_/A VGND VGND VPWR VPWR _10586_/Y sky130_fd_sc_hd__inv_2
X_16093_ _16031_/X _16092_/Y _16031_/X _16092_/Y VGND VGND VPWR VPWR _16213_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12256_ _12256_/A _12256_/B VGND VGND VPWR VPWR _12256_/Y sky130_fd_sc_hd__nor2_1
X_15044_ _15044_/A _15044_/B VGND VGND VPWR VPWR _15044_/X sky130_fd_sc_hd__or2_1
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11207_ _11207_/A _11220_/B VGND VGND VPWR VPWR _13331_/A sky130_fd_sc_hd__or2_1
X_12187_ _13712_/A _12261_/B _12261_/A _12261_/B VGND VGND VPWR VPWR _12187_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11138_ _11138_/A _12089_/A VGND VGND VPWR VPWR _11138_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15946_ _14370_/X _14372_/Y _15839_/B _14374_/A _14369_/A VGND VGND VPWR VPWR _15947_/B
+ sky130_fd_sc_hd__o221a_1
X_11069_ _12827_/A VGND VGND VPWR VPWR _12915_/A sky130_fd_sc_hd__buf_1
X_15877_ _15890_/A _15890_/B VGND VGND VPWR VPWR _15877_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14828_ _15437_/A VGND VGND VPWR VPWR _14930_/A sky130_fd_sc_hd__buf_1
XFILLER_63_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14759_ _14750_/X _14758_/X _14750_/X _14758_/X VGND VGND VPWR VPWR _14761_/B sky130_fd_sc_hd__a2bb2o_1
X_08280_ input2/X VGND VGND VPWR VPWR _08358_/A sky130_fd_sc_hd__inv_4
X_16429_ _16447_/A _16429_/B VGND VGND VPWR VPWR _16429_/X sky130_fd_sc_hd__or2_1
XFILLER_32_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09803_ _09803_/A _09803_/B VGND VGND VPWR VPWR _09856_/B sky130_fd_sc_hd__or2_1
XFILLER_75_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09734_ _09734_/A _09734_/B VGND VGND VPWR VPWR _09737_/B sky130_fd_sc_hd__or2_1
XFILLER_67_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09665_ _09579_/Y _09663_/X _09664_/Y VGND VGND VPWR VPWR _09665_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08616_ _09221_/A VGND VGND VPWR VPWR _08716_/A sky130_fd_sc_hd__inv_2
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09596_ _09554_/X _09595_/Y _09554_/X _09595_/Y VGND VGND VPWR VPWR _09658_/B sky130_fd_sc_hd__a2bb2o_1
X_08547_ _08546_/A _08446_/Y _08546_/Y _08446_/A VGND VGND VPWR VPWR _10118_/B sky130_fd_sc_hd__o22a_1
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08478_ input28/X input12/X VGND VGND VPWR VPWR _08478_/Y sky130_fd_sc_hd__nor2_1
X_10440_ _10440_/A VGND VGND VPWR VPWR _11848_/A sky130_fd_sc_hd__buf_1
XFILLER_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10371_ _09415_/A _09118_/B _09118_/Y VGND VGND VPWR VPWR _10371_/X sky130_fd_sc_hd__o21a_1
X_12110_ _13198_/A _12065_/B _12065_/Y VGND VGND VPWR VPWR _12110_/Y sky130_fd_sc_hd__o21ai_1
X_13090_ _13090_/A _13015_/X VGND VGND VPWR VPWR _13090_/X sky130_fd_sc_hd__or2b_1
XFILLER_123_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12041_ _11965_/X _12040_/X _11965_/X _12040_/X VGND VGND VPWR VPWR _12051_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15800_ _16099_/A _15800_/B VGND VGND VPWR VPWR _15800_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13992_ _13989_/X _13991_/X _13989_/X _13991_/X VGND VGND VPWR VPWR _13994_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15731_ _16114_/A _15815_/B VGND VGND VPWR VPWR _15731_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12943_ _12880_/Y _12941_/X _12942_/Y VGND VGND VPWR VPWR _12943_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15662_ _15947_/A _15662_/B VGND VGND VPWR VPWR _15662_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12874_ _12857_/A _12857_/B _12857_/Y VGND VGND VPWR VPWR _12874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15593_ _15503_/X _15593_/B VGND VGND VPWR VPWR _15593_/X sky130_fd_sc_hd__and2b_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _15345_/A _14659_/B VGND VGND VPWR VPWR _14613_/Y sky130_fd_sc_hd__nor2_1
X_11825_ _10396_/A _11778_/B _10396_/A _11778_/B VGND VGND VPWR VPWR _11825_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14544_/A _14519_/X VGND VGND VPWR VPWR _14544_/X sky130_fd_sc_hd__or2b_1
XFILLER_60_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11756_ _11775_/B VGND VGND VPWR VPWR _11756_/Y sky130_fd_sc_hd__inv_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _14470_/X _14474_/X _14470_/X _14474_/X VGND VGND VPWR VPWR _14476_/B sky130_fd_sc_hd__a2bb2o_1
X_10707_ _10785_/A _10706_/Y _10785_/A _10706_/Y VGND VGND VPWR VPWR _10708_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16214_ _16214_/A VGND VGND VPWR VPWR _16214_/Y sky130_fd_sc_hd__inv_2
X_13426_ _13422_/Y _13424_/Y _13425_/Y VGND VGND VPWR VPWR _13430_/B sky130_fd_sc_hd__o21ai_1
X_11687_ _12431_/A _11626_/A _11627_/Y _11630_/X VGND VGND VPWR VPWR _11687_/X sky130_fd_sc_hd__o22a_1
XFILLER_127_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10638_ _11882_/A VGND VGND VPWR VPWR _12992_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16145_ _16273_/A _16272_/A VGND VGND VPWR VPWR _16145_/Y sky130_fd_sc_hd__nor2_1
X_13357_ _15467_/A _13344_/B _13344_/Y _13356_/X VGND VGND VPWR VPWR _13357_/X sky130_fd_sc_hd__o2bb2a_1
X_10569_ _10557_/X _10568_/Y _10557_/X _10568_/Y VGND VGND VPWR VPWR _10675_/A sky130_fd_sc_hd__o2bb2a_1
X_16076_ _16108_/A _16108_/B VGND VGND VPWR VPWR _16076_/X sky130_fd_sc_hd__and2_1
X_12308_ _12308_/A _12308_/B VGND VGND VPWR VPWR _12308_/Y sky130_fd_sc_hd__nand2_1
X_13288_ _14732_/A _13288_/B VGND VGND VPWR VPWR _13288_/Y sky130_fd_sc_hd__nand2_1
X_12239_ _13350_/A _12238_/B _12237_/X _12238_/Y VGND VGND VPWR VPWR _12239_/X sky130_fd_sc_hd__a2bb2o_1
X_15027_ _12830_/A _12830_/B _10426_/A _12830_/Y VGND VGND VPWR VPWR _15027_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 wbs_adr_i[11] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_8
X_15929_ _15895_/X _15928_/Y _15895_/X _15928_/Y VGND VGND VPWR VPWR _15958_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09450_ _09484_/A _09527_/A VGND VGND VPWR VPWR _09450_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08401_ _08401_/A _09677_/B VGND VGND VPWR VPWR _08670_/A sky130_fd_sc_hd__or2_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09381_ _10240_/A VGND VGND VPWR VPWR _09382_/B sky130_fd_sc_hd__buf_1
X_08332_ _08332_/A _08332_/B VGND VGND VPWR VPWR _08333_/A sky130_fd_sc_hd__or2_1
X_08263_ _08263_/A input14/X VGND VGND VPWR VPWR _08342_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09717_ _09717_/A _09717_/B VGND VGND VPWR VPWR _09717_/X sky130_fd_sc_hd__or2_1
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09648_ _09648_/A _09648_/B VGND VGND VPWR VPWR _09648_/Y sky130_fd_sc_hd__nor2_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09579_ _09995_/A _09664_/B VGND VGND VPWR VPWR _09579_/Y sky130_fd_sc_hd__nor2_1
X_12590_ _12590_/A VGND VGND VPWR VPWR _12590_/Y sky130_fd_sc_hd__inv_2
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11610_/A VGND VGND VPWR VPWR _11610_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11541_ _13495_/A _11629_/B _13495_/A _11629_/B VGND VGND VPWR VPWR _11541_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14260_ _14215_/Y _14258_/Y _14259_/Y VGND VGND VPWR VPWR _14261_/A sky130_fd_sc_hd__o21ai_2
XFILLER_109_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11472_ _13313_/A VGND VGND VPWR VPWR _14005_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14191_ _15860_/A _14271_/B VGND VGND VPWR VPWR _14191_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13211_ _15107_/A VGND VGND VPWR VPWR _14841_/A sky130_fd_sc_hd__inv_2
X_10423_ _10423_/A VGND VGND VPWR VPWR _10424_/B sky130_fd_sc_hd__inv_2
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13142_ _14953_/A _13125_/B _13125_/Y VGND VGND VPWR VPWR _13142_/Y sky130_fd_sc_hd__o21ai_1
X_10354_ _10424_/A _10421_/B VGND VGND VPWR VPWR _10354_/X sky130_fd_sc_hd__or2_1
XFILLER_112_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13073_ _13073_/A VGND VGND VPWR VPWR _13764_/A sky130_fd_sc_hd__inv_2
X_10285_ _10282_/A _10281_/A _10350_/A _10284_/Y VGND VGND VPWR VPWR _10286_/B sky130_fd_sc_hd__o22a_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12024_ _13194_/A _12061_/B VGND VGND VPWR VPWR _12024_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13975_ _13865_/X _13974_/Y _13875_/Y VGND VGND VPWR VPWR _13997_/A sky130_fd_sc_hd__o21ai_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15714_ _14925_/X _15713_/X _14925_/X _15713_/X VGND VGND VPWR VPWR _15715_/B sky130_fd_sc_hd__a2bb2oi_1
X_12926_ _14458_/A _12926_/B VGND VGND VPWR VPWR _12926_/Y sky130_fd_sc_hd__nand2_1
X_15645_ _14378_/X _15644_/Y _14378_/X _15644_/Y VGND VGND VPWR VPWR _15669_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12857_ _12857_/A _12857_/B VGND VGND VPWR VPWR _12857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11808_ _11808_/A _11808_/B VGND VGND VPWR VPWR _11808_/Y sky130_fd_sc_hd__nor2_1
X_15576_ _15972_/A _14402_/B _14402_/Y VGND VGND VPWR VPWR _15576_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _12724_/Y _12787_/X _12724_/Y _12787_/X VGND VGND VPWR VPWR _12789_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14527_ _12003_/Y _14526_/X _12003_/Y _14526_/X VGND VGND VPWR VPWR _14528_/B sky130_fd_sc_hd__o2bb2a_1
X_11739_ _11745_/A _11746_/A VGND VGND VPWR VPWR _11739_/Y sky130_fd_sc_hd__nor2_1
X_14458_ _14458_/A _14458_/B VGND VGND VPWR VPWR _14458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14389_ _15960_/A _14389_/B VGND VGND VPWR VPWR _15605_/B sky130_fd_sc_hd__or2_1
X_13409_ _13355_/Y _13408_/X _13355_/Y _13408_/X VGND VGND VPWR VPWR _13410_/A sky130_fd_sc_hd__a2bb2o_1
X_16128_ _16126_/Y _16127_/X _16126_/Y _16127_/X VGND VGND VPWR VPWR _16128_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_115_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16059_ _15995_/X _16059_/B VGND VGND VPWR VPWR _16059_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08950_ _09539_/A _08647_/A _08648_/X VGND VGND VPWR VPWR _08950_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08881_ _08881_/A _08881_/B VGND VGND VPWR VPWR _08881_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09502_ _09502_/A _09502_/B VGND VGND VPWR VPWR _09502_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09433_ _09766_/A _09433_/B VGND VGND VPWR VPWR _09433_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _09429_/B _11577_/A VGND VGND VPWR VPWR _09364_/X sky130_fd_sc_hd__or2_1
XFILLER_52_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08315_ _08313_/Y _08314_/A _08313_/A _08314_/Y _08304_/X VGND VGND VPWR VPWR _08532_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09295_ _09629_/A _09294_/X _09629_/A _09294_/X VGND VGND VPWR VPWR _09296_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08246_ input4/X VGND VGND VPWR VPWR _08316_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10070_ _10022_/X _10069_/Y _10022_/X _10069_/Y VGND VGND VPWR VPWR _10071_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13760_ _13760_/A _13760_/B VGND VGND VPWR VPWR _13760_/X sky130_fd_sc_hd__or2_1
X_10972_ _10972_/A VGND VGND VPWR VPWR _12176_/A sky130_fd_sc_hd__inv_2
XFILLER_16_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13691_ _13672_/Y _13689_/X _13690_/Y VGND VGND VPWR VPWR _13691_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12711_ _12704_/A _12704_/B _12704_/X _12710_/X VGND VGND VPWR VPWR _12711_/X sky130_fd_sc_hd__o22a_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12642_ _12642_/A VGND VGND VPWR VPWR _12642_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15430_ _14971_/A _15167_/B _15167_/Y _15169_/Y VGND VGND VPWR VPWR _15430_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12573_ _12573_/A VGND VGND VPWR VPWR _12573_/Y sky130_fd_sc_hd__inv_2
X_15361_ _15350_/X _15360_/Y _15350_/X _15360_/Y VGND VGND VPWR VPWR _15418_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14312_ _13439_/A _13439_/B _13439_/Y VGND VGND VPWR VPWR _14312_/X sky130_fd_sc_hd__o21a_1
X_15292_ _15283_/X _15291_/Y _15283_/X _15291_/Y VGND VGND VPWR VPWR _15353_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11524_ _10086_/X _11523_/X _10086_/X _11523_/X VGND VGND VPWR VPWR _11525_/B sky130_fd_sc_hd__a2bb2o_1
X_14243_ _14243_/A _14243_/B VGND VGND VPWR VPWR _14361_/B sky130_fd_sc_hd__or2_1
X_11455_ _15540_/A _11455_/B VGND VGND VPWR VPWR _11455_/Y sky130_fd_sc_hd__nand2_1
X_10406_ _11783_/A VGND VGND VPWR VPWR _13567_/A sky130_fd_sc_hd__buf_1
XFILLER_125_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14174_ _14127_/X _14173_/Y _14127_/X _14173_/Y VGND VGND VPWR VPWR _14175_/B sky130_fd_sc_hd__a2bb2oi_1
X_11386_ _12314_/A _11386_/B VGND VGND VPWR VPWR _11386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13125_ _15234_/A _13125_/B VGND VGND VPWR VPWR _13125_/Y sky130_fd_sc_hd__nand2_1
X_10337_ _10291_/B _10336_/Y _10291_/B _10336_/Y VGND VGND VPWR VPWR _10338_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13056_ _13028_/X _13055_/X _13028_/X _13055_/X VGND VGND VPWR VPWR _13119_/B sky130_fd_sc_hd__a2bb2o_1
X_10268_ _10268_/A VGND VGND VPWR VPWR _10471_/A sky130_fd_sc_hd__clkbuf_2
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12007_ _12007_/A _12073_/B VGND VGND VPWR VPWR _12007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10199_ _10196_/X _10198_/X _10196_/X _10198_/X VGND VGND VPWR VPWR _10346_/B sky130_fd_sc_hd__o2bb2a_4
X_13958_ _13896_/Y _13956_/X _13957_/Y VGND VGND VPWR VPWR _13958_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12909_ _13608_/A VGND VGND VPWR VPWR _12925_/A sky130_fd_sc_hd__buf_1
XFILLER_46_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13889_ _13889_/A VGND VGND VPWR VPWR _15418_/A sky130_fd_sc_hd__buf_1
XFILLER_62_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _14341_/X _15628_/B VGND VGND VPWR VPWR _15628_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15559_ _15430_/X _15558_/X _15430_/X _15558_/X VGND VGND VPWR VPWR _15559_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09080_ _09760_/A VGND VGND VPWR VPWR _09432_/A sky130_fd_sc_hd__buf_1
XFILLER_128_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09982_ _09700_/Y _09980_/Y _09981_/Y VGND VGND VPWR VPWR _09984_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08933_ _10228_/B _08932_/B _08931_/Y _08932_/Y VGND VGND VPWR VPWR _08942_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08864_ _09490_/A _08792_/Y _08793_/Y _08863_/X VGND VGND VPWR VPWR _08864_/X sky130_fd_sc_hd__o22a_1
X_08795_ _09492_/A VGND VGND VPWR VPWR _08795_/X sky130_fd_sc_hd__buf_1
XFILLER_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09416_ _09946_/A _09414_/Y _09415_/Y VGND VGND VPWR VPWR _09418_/B sky130_fd_sc_hd__o21ai_1
XFILLER_13_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09347_ _09525_/A _09347_/B VGND VGND VPWR VPWR _09348_/A sky130_fd_sc_hd__or2_1
X_09278_ _10254_/A VGND VGND VPWR VPWR _09312_/A sky130_fd_sc_hd__buf_1
X_08229_ _08229_/A VGND VGND VPWR VPWR _08230_/A sky130_fd_sc_hd__buf_1
XFILLER_126_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11240_ _14042_/A VGND VGND VPWR VPWR _12232_/A sky130_fd_sc_hd__inv_2
XFILLER_4_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11171_ _12195_/A _11170_/B _11170_/Y VGND VGND VPWR VPWR _11171_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10122_ _10237_/B VGND VGND VPWR VPWR _10122_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14930_ _14930_/A _14930_/B VGND VGND VPWR VPWR _14930_/X sky130_fd_sc_hd__and2_1
XFILLER_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10053_ _09066_/A _09681_/A _09401_/Y _08931_/A VGND VGND VPWR VPWR _10055_/A sky130_fd_sc_hd__o22a_1
X_14861_ _14930_/A _14930_/B _14930_/A _14930_/B VGND VGND VPWR VPWR _14861_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13812_ _13812_/A _13766_/X VGND VGND VPWR VPWR _13812_/X sky130_fd_sc_hd__or2b_1
XFILLER_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14792_ _14792_/A _14732_/X VGND VGND VPWR VPWR _14792_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13743_ _13760_/A _13760_/B VGND VGND VPWR VPWR _13821_/A sky130_fd_sc_hd__and2_1
XFILLER_73_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10955_ _11990_/A _10955_/B VGND VGND VPWR VPWR _10955_/X sky130_fd_sc_hd__and2_1
XFILLER_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16462_ _16357_/A _16462_/D VGND VGND VPWR VPWR _16462_/Q sky130_fd_sc_hd__dfxtp_1
X_10886_ _10886_/A _10886_/B VGND VGND VPWR VPWR _10886_/X sky130_fd_sc_hd__and2_1
X_13674_ _13618_/X _13673_/X _13618_/X _13673_/X VGND VGND VPWR VPWR _13688_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16393_ _16402_/A VGND VGND VPWR VPWR _16393_/Y sky130_fd_sc_hd__inv_2
X_12625_ _14213_/A _12623_/X _12624_/X VGND VGND VPWR VPWR _12625_/X sky130_fd_sc_hd__o21a_1
X_15413_ _15447_/A _15411_/X _15412_/X VGND VGND VPWR VPWR _15413_/X sky130_fd_sc_hd__o21a_1
X_12556_ _12556_/A VGND VGND VPWR VPWR _12556_/Y sky130_fd_sc_hd__inv_2
X_15344_ _15372_/A _15342_/X _15343_/X VGND VGND VPWR VPWR _15344_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11507_ _11506_/A _11506_/B _11506_/X _11305_/X VGND VGND VPWR VPWR _11635_/A sky130_fd_sc_hd__o22a_1
XFILLER_8_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12487_ _14065_/A _12407_/B _12407_/Y _12358_/X VGND VGND VPWR VPWR _12487_/Y sky130_fd_sc_hd__a2bb2oi_1
X_15275_ _14577_/A _15261_/B _15261_/Y _15274_/X VGND VGND VPWR VPWR _15275_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14226_ _12619_/X _14225_/Y _12619_/X _14225_/Y VGND VGND VPWR VPWR _14253_/B sky130_fd_sc_hd__a2bb2o_1
X_11438_ _11433_/Y _12576_/A _11437_/Y VGND VGND VPWR VPWR _11443_/B sky130_fd_sc_hd__o21ai_1
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14157_ _14230_/A VGND VGND VPWR VPWR _14206_/A sky130_fd_sc_hd__clkbuf_2
X_11369_ _12308_/A VGND VGND VPWR VPWR _14125_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13108_ _13087_/Y _13106_/X _13107_/Y VGND VGND VPWR VPWR _13108_/X sky130_fd_sc_hd__o21a_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14088_ _13344_/A _14038_/B _14038_/A _14038_/B VGND VGND VPWR VPWR _14088_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13039_ _13882_/A VGND VGND VPWR VPWR _15234_/A sky130_fd_sc_hd__buf_1
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08580_ _09323_/A _09209_/B _10013_/A _08579_/Y VGND VGND VPWR VPWR _08580_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09201_ _09193_/Y _09200_/X _09193_/Y _09200_/X VGND VGND VPWR VPWR _11413_/B sky130_fd_sc_hd__a2bb2o_4
X_09132_ _09128_/Y _09130_/Y _09131_/Y VGND VGND VPWR VPWR _09136_/B sky130_fd_sc_hd__o21ai_1
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09063_ _08839_/A _09042_/X _08839_/A _09042_/X VGND VGND VPWR VPWR _09070_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09965_ _09995_/A _09995_/B VGND VGND VPWR VPWR _09965_/X sky130_fd_sc_hd__and2_1
XFILLER_134_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _09882_/A _09882_/B _09883_/B VGND VGND VPWR VPWR _09898_/A sky130_fd_sc_hd__a21bo_1
X_08916_ _08916_/A _09817_/B VGND VGND VPWR VPWR _08917_/A sky130_fd_sc_hd__or2_1
XFILLER_97_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _08847_/A VGND VGND VPWR VPWR _09503_/B sky130_fd_sc_hd__buf_1
XFILLER_18_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08778_ _08778_/A _10131_/A VGND VGND VPWR VPWR _08778_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10740_ _10637_/A _10739_/Y _10637_/A _10739_/Y VGND VGND VPWR VPWR _10741_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10671_ _10077_/A _10670_/Y _09969_/Y _10670_/A _10959_/A VGND VGND VPWR VPWR _11919_/A
+ sky130_fd_sc_hd__o221a_1
X_12410_ _12410_/A _12410_/B VGND VGND VPWR VPWR _12410_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13390_ _13390_/A _13362_/X VGND VGND VPWR VPWR _13390_/X sky130_fd_sc_hd__or2b_1
X_12341_ _13395_/A _12341_/B VGND VGND VPWR VPWR _12341_/Y sky130_fd_sc_hd__nand2_1
X_15060_ _15060_/A _15060_/B VGND VGND VPWR VPWR _15060_/Y sky130_fd_sc_hd__nand2_1
X_12272_ _12272_/A VGND VGND VPWR VPWR _12272_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14011_ _14011_/A _14061_/B VGND VGND VPWR VPWR _14011_/X sky130_fd_sc_hd__and2_1
X_11223_ _11223_/A _11084_/X VGND VGND VPWR VPWR _11223_/X sky130_fd_sc_hd__or2b_1
XFILLER_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11154_ _09382_/B _10240_/B _10240_/X VGND VGND VPWR VPWR _11155_/B sky130_fd_sc_hd__a21boi_1
XFILLER_122_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15962_ _15962_/A _15962_/B VGND VGND VPWR VPWR _16002_/B sky130_fd_sc_hd__or2_1
XFILLER_110_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11085_ _11223_/A _11083_/X _11084_/X VGND VGND VPWR VPWR _11085_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10105_ _08671_/A _10105_/A2 _09627_/A _08667_/Y VGND VGND VPWR VPWR _10177_/B sky130_fd_sc_hd__o22a_1
X_14913_ _14892_/Y _14911_/X _14912_/Y VGND VGND VPWR VPWR _14913_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10036_ _10029_/X _10035_/Y _10029_/X _10035_/Y VGND VGND VPWR VPWR _10087_/B sky130_fd_sc_hd__a2bb2o_1
X_15893_ _15874_/Y _15891_/X _15892_/Y VGND VGND VPWR VPWR _15893_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14844_ _14944_/A _14944_/B VGND VGND VPWR VPWR _14844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14775_ _15443_/A VGND VGND VPWR VPWR _14778_/A sky130_fd_sc_hd__buf_1
X_11987_ _11987_/A _11987_/B VGND VGND VPWR VPWR _11987_/X sky130_fd_sc_hd__or2_1
XFILLER_17_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13726_ _13726_/A _13700_/X VGND VGND VPWR VPWR _13726_/X sky130_fd_sc_hd__or2b_1
X_10938_ _12070_/A _10938_/B VGND VGND VPWR VPWR _10938_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16445_ _16445_/A _16445_/B VGND VGND VPWR VPWR _16445_/X sky130_fd_sc_hd__and2_1
X_10869_ _10776_/X _10868_/Y _10776_/X _10868_/Y VGND VGND VPWR VPWR _10870_/B sky130_fd_sc_hd__o2bb2a_1
X_13657_ _13700_/A _13700_/B VGND VGND VPWR VPWR _13726_/A sky130_fd_sc_hd__and2_1
X_16376_ _16319_/X _16375_/Y _16319_/X _16375_/Y VGND VGND VPWR VPWR _16397_/A sky130_fd_sc_hd__a2bb2o_1
X_12608_ _14243_/A _12608_/B VGND VGND VPWR VPWR _12608_/Y sky130_fd_sc_hd__nand2_1
X_13588_ _13579_/X _13587_/Y _13579_/X _13587_/Y VGND VGND VPWR VPWR _13637_/B sky130_fd_sc_hd__a2bb2o_1
X_12539_ _13437_/A _11386_/B _11386_/Y VGND VGND VPWR VPWR _12540_/B sky130_fd_sc_hd__o21a_1
X_15327_ _14567_/A _15270_/B _14567_/A _15270_/B VGND VGND VPWR VPWR _15327_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15258_ _15258_/A _15258_/B VGND VGND VPWR VPWR _15258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14209_ _15869_/A _14262_/B VGND VGND VPWR VPWR _14209_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15189_ _15154_/X _15188_/Y _15154_/X _15188_/Y VGND VGND VPWR VPWR _15190_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09750_ _09750_/A _09750_/B VGND VGND VPWR VPWR _09750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ _08701_/A _08701_/B VGND VGND VPWR VPWR _08703_/A sky130_fd_sc_hd__or2_2
X_09681_ _09681_/A _09681_/B VGND VGND VPWR VPWR _09684_/B sky130_fd_sc_hd__or2_1
XFILLER_104_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08632_ _09251_/A _09225_/B _10017_/A _08631_/Y VGND VGND VPWR VPWR _08632_/X sky130_fd_sc_hd__o22a_1
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08563_ _08589_/A _08563_/B VGND VGND VPWR VPWR _09453_/B sky130_fd_sc_hd__or2_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08494_ _08311_/A _08245_/B _08470_/Y _08516_/A VGND VGND VPWR VPWR _08501_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09115_ _09415_/A _09118_/B VGND VGND VPWR VPWR _09115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09046_ _08715_/A _08715_/B _08715_/X _09045_/X VGND VGND VPWR VPWR _09047_/A sky130_fd_sc_hd__a22o_1
XFILLER_123_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09948_ _09946_/A _09947_/A _09946_/Y _09947_/Y _09391_/A VGND VGND VPWR VPWR _09949_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09879_ _09867_/X _08789_/Y _09867_/X _08789_/Y VGND VGND VPWR VPWR _09884_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11910_ _11910_/A _11910_/B VGND VGND VPWR VPWR _11910_/Y sky130_fd_sc_hd__nand2_1
X_12890_ _12849_/A _12849_/B _12849_/Y VGND VGND VPWR VPWR _12890_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11841_ _11830_/Y _11839_/X _11840_/Y VGND VGND VPWR VPWR _11841_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _14560_/A _14511_/X VGND VGND VPWR VPWR _14560_/X sky130_fd_sc_hd__or2b_1
XFILLER_54_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11772_ _11801_/B _11771_/Y _11801_/B _11771_/Y VGND VGND VPWR VPWR _11773_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10644_/A _10722_/Y _10644_/A _10722_/Y VGND VGND VPWR VPWR _10724_/B sky130_fd_sc_hd__a2bb2o_1
X_13511_ _10696_/X _13486_/X _10696_/X _13486_/X VGND VGND VPWR VPWR _13512_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14491_ _15202_/A _14515_/B VGND VGND VPWR VPWR _14552_/A sky130_fd_sc_hd__and2_1
XFILLER_41_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16230_ _16251_/B VGND VGND VPWR VPWR _16318_/A sky130_fd_sc_hd__clkbuf_2
X_13442_ _13386_/Y _13440_/X _13441_/Y VGND VGND VPWR VPWR _13442_/X sky130_fd_sc_hd__o21a_1
X_10654_ _13632_/A _10654_/B VGND VGND VPWR VPWR _10654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16161_ _16268_/B VGND VGND VPWR VPWR _16334_/A sky130_fd_sc_hd__buf_6
X_13373_ _13310_/X _13372_/X _13310_/X _13372_/X VGND VGND VPWR VPWR _13449_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10585_ _09723_/A _09723_/B _09723_/Y VGND VGND VPWR VPWR _10586_/A sky130_fd_sc_hd__o21ai_1
X_12324_ _12324_/A _12324_/B VGND VGND VPWR VPWR _12324_/X sky130_fd_sc_hd__and2_1
X_15112_ _15098_/X _15111_/Y _15098_/X _15111_/Y VGND VGND VPWR VPWR _15113_/B sky130_fd_sc_hd__a2bb2o_1
X_16092_ _16032_/A _16032_/B _16032_/Y VGND VGND VPWR VPWR _16092_/Y sky130_fd_sc_hd__o21ai_1
X_12255_ _12254_/Y _12161_/X _12195_/Y VGND VGND VPWR VPWR _12255_/X sky130_fd_sc_hd__o21a_1
X_15043_ _15061_/A _15041_/X _15042_/X VGND VGND VPWR VPWR _15043_/X sky130_fd_sc_hd__o21a_1
X_11206_ _14055_/A _11206_/B VGND VGND VPWR VPWR _11206_/Y sky130_fd_sc_hd__nand2_1
X_12186_ _12263_/B _12185_/Y _12263_/B _12185_/Y VGND VGND VPWR VPWR _12261_/B sky130_fd_sc_hd__o2bb2a_1
X_11137_ _12174_/A VGND VGND VPWR VPWR _12089_/A sky130_fd_sc_hd__inv_2
XFILLER_1_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15945_ _15948_/A _15948_/B VGND VGND VPWR VPWR _15945_/X sky130_fd_sc_hd__and2_1
X_11068_ _11246_/A VGND VGND VPWR VPWR _12234_/B sky130_fd_sc_hd__inv_2
XFILLER_76_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15876_ _14219_/X _15842_/X _14219_/X _15842_/X VGND VGND VPWR VPWR _15890_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10019_ _08935_/A _09069_/A _08917_/A _08935_/X VGND VGND VPWR VPWR _10019_/X sky130_fd_sc_hd__a22o_1
X_14827_ _14774_/A _14774_/B _14774_/X _14826_/X VGND VGND VPWR VPWR _14827_/X sky130_fd_sc_hd__o22a_1
XFILLER_91_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14758_ _14757_/A _14757_/B _14757_/Y VGND VGND VPWR VPWR _14758_/X sky130_fd_sc_hd__a21o_1
X_14689_ _14740_/A _14740_/B VGND VGND VPWR VPWR _14776_/A sky130_fd_sc_hd__and2_1
X_13709_ _12855_/A _13648_/B _13708_/Y _13645_/X VGND VGND VPWR VPWR _13709_/X sky130_fd_sc_hd__o22a_1
X_16428_ _16470_/Q VGND VGND VPWR VPWR _16428_/Y sky130_fd_sc_hd__inv_2
X_16359_ _16330_/A _16330_/B _16330_/Y VGND VGND VPWR VPWR _16359_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09802_ _09802_/A _09844_/A VGND VGND VPWR VPWR _09803_/B sky130_fd_sc_hd__or2_1
XFILLER_101_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09733_ _09733_/A _09733_/B VGND VGND VPWR VPWR _09736_/A sky130_fd_sc_hd__or2_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09664_ _09995_/A _09664_/B VGND VGND VPWR VPWR _09664_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08615_ _09457_/B VGND VGND VPWR VPWR _09547_/A sky130_fd_sc_hd__buf_1
X_09595_ _09595_/A _09595_/B VGND VGND VPWR VPWR _09595_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08546_ _08546_/A VGND VGND VPWR VPWR _08546_/Y sky130_fd_sc_hd__inv_2
X_08477_ input29/X input13/X VGND VGND VPWR VPWR _08477_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10370_ _10369_/Y _10309_/Y _10307_/Y VGND VGND VPWR VPWR _10370_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09029_ _09029_/A _09540_/B VGND VGND VPWR VPWR _09030_/B sky130_fd_sc_hd__or2_1
X_12040_ _12040_/A _11966_/X VGND VGND VPWR VPWR _12040_/X sky130_fd_sc_hd__or2b_1
XFILLER_78_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13991_ _13860_/X _13990_/Y _13885_/Y VGND VGND VPWR VPWR _13991_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15730_ _15682_/X _15729_/Y _15682_/X _15729_/Y VGND VGND VPWR VPWR _15815_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12942_ _12942_/A _12942_/B VGND VGND VPWR VPWR _12942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15661_ _15661_/A VGND VGND VPWR VPWR _15947_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14612_ _14586_/X _14611_/Y _14586_/X _14611_/Y VGND VGND VPWR VPWR _14659_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12873_ _12944_/A VGND VGND VPWR VPWR _14676_/A sky130_fd_sc_hd__buf_1
XFILLER_61_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15592_ _15683_/A _15683_/B VGND VGND VPWR VPWR _15592_/Y sky130_fd_sc_hd__nor2_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11824_ _13624_/A _11844_/B VGND VGND VPWR VPWR _11824_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14543_ _15252_/A VGND VGND VPWR VPWR _14583_/A sky130_fd_sc_hd__buf_1
X_11755_ _11760_/B _11754_/Y _11760_/B _11754_/Y VGND VGND VPWR VPWR _11775_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14474_ _14473_/A _14473_/B _14473_/Y VGND VGND VPWR VPWR _14474_/X sky130_fd_sc_hd__a21o_1
X_10706_ _13698_/A _10784_/B _10705_/Y VGND VGND VPWR VPWR _10706_/Y sky130_fd_sc_hd__o21ai_1
X_16213_ _16213_/A VGND VGND VPWR VPWR _16213_/Y sky130_fd_sc_hd__inv_2
X_13425_ _14100_/A _13425_/B VGND VGND VPWR VPWR _13425_/Y sky130_fd_sc_hd__nand2_1
X_11686_ _15163_/A VGND VGND VPWR VPWR _12431_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10637_ _10637_/A VGND VGND VPWR VPWR _10637_/Y sky130_fd_sc_hd__inv_2
X_16144_ _16160_/A _16144_/B VGND VGND VPWR VPWR _16272_/A sky130_fd_sc_hd__or2_1
X_13356_ _15470_/A _13348_/B _13348_/Y _13355_/Y VGND VGND VPWR VPWR _13356_/X sky130_fd_sc_hd__o2bb2a_1
X_10568_ _10568_/A VGND VGND VPWR VPWR _10568_/Y sky130_fd_sc_hd__clkinvlp_2
X_16075_ _16039_/X _16074_/Y _16039_/X _16074_/Y VGND VGND VPWR VPWR _16108_/B sky130_fd_sc_hd__a2bb2o_1
X_12307_ _12247_/X _12306_/Y _12247_/X _12306_/Y VGND VGND VPWR VPWR _12308_/B sky130_fd_sc_hd__a2bb2o_1
X_13287_ _13287_/A VGND VGND VPWR VPWR _13287_/Y sky130_fd_sc_hd__inv_2
X_10499_ _10499_/A VGND VGND VPWR VPWR _10499_/Y sky130_fd_sc_hd__inv_2
X_12238_ _13350_/A _12238_/B VGND VGND VPWR VPWR _12238_/Y sky130_fd_sc_hd__nand2_1
X_15026_ _15028_/A _15028_/B VGND VGND VPWR VPWR _15082_/A sky130_fd_sc_hd__and2_1
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12169_ _12169_/A _12169_/B VGND VGND VPWR VPWR _12169_/X sky130_fd_sc_hd__or2_1
XFILLER_84_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15928_ _15896_/A _15896_/B _15896_/Y VGND VGND VPWR VPWR _15928_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 wbs_adr_i[12] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_2
XFILLER_37_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15859_ _15902_/A _15902_/B VGND VGND VPWR VPWR _15859_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08400_ _08662_/B _08400_/B VGND VGND VPWR VPWR _09677_/B sky130_fd_sc_hd__or2_1
X_09380_ _09334_/X _08883_/Y _09334_/X _08883_/Y VGND VGND VPWR VPWR _10240_/A sky130_fd_sc_hd__o2bb2a_1
X_08331_ _08331_/A input32/X VGND VGND VPWR VPWR _08332_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08262_ input30/X VGND VGND VPWR VPWR _08263_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_20_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09716_ _09716_/A _09717_/B VGND VGND VPWR VPWR _10597_/A sky130_fd_sc_hd__and2_1
XFILLER_28_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09647_ _09975_/A _09650_/B VGND VGND VPWR VPWR _09647_/Y sky130_fd_sc_hd__nor2_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09558_/X _09577_/X _09558_/X _09577_/X VGND VGND VPWR VPWR _09664_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08701_/A _08529_/B VGND VGND VPWR VPWR _09527_/A sky130_fd_sc_hd__or2_2
X_11540_ _11520_/X _11539_/X _11520_/X _11539_/X VGND VGND VPWR VPWR _11629_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11471_ _09184_/Y _11470_/A _09184_/A _11470_/Y _09204_/X VGND VGND VPWR VPWR _13313_/A
+ sky130_fd_sc_hd__a221o_4
X_14190_ _12631_/X _14189_/X _12631_/X _14189_/X VGND VGND VPWR VPWR _14271_/B sky130_fd_sc_hd__a2bb2o_1
X_13210_ _14934_/A _13451_/B _13209_/Y VGND VGND VPWR VPWR _13210_/Y sky130_fd_sc_hd__o21ai_1
X_10422_ _10422_/A VGND VGND VPWR VPWR _10426_/A sky130_fd_sc_hd__inv_2
XFILLER_109_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13141_ _15234_/A VGND VGND VPWR VPWR _14953_/A sky130_fd_sc_hd__buf_1
X_10353_ _10423_/A VGND VGND VPWR VPWR _10421_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13072_ _15252_/A _13113_/B VGND VGND VPWR VPWR _13072_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12023_ _11975_/X _12022_/Y _11975_/X _12022_/Y VGND VGND VPWR VPWR _12061_/B sky130_fd_sc_hd__a2bb2o_1
X_10284_ _13478_/B VGND VGND VPWR VPWR _10284_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15713_ _15550_/A _14926_/B _14926_/Y VGND VGND VPWR VPWR _15713_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13974_ _13974_/A _13974_/B VGND VGND VPWR VPWR _13974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12925_ _12925_/A VGND VGND VPWR VPWR _14458_/A sky130_fd_sc_hd__buf_1
XFILLER_34_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15644_ _14353_/X _15644_/B VGND VGND VPWR VPWR _15644_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_61_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12856_ _12802_/Y _12854_/X _12855_/Y VGND VGND VPWR VPWR _12856_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15575_ _15700_/A _15575_/B VGND VGND VPWR VPWR _16055_/A sky130_fd_sc_hd__or2_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11806_/A _11806_/B _11806_/X _11767_/B VGND VGND VPWR VPWR _11855_/B sky130_fd_sc_hd__a22o_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _15040_/A _11988_/Y _11931_/Y _14471_/X VGND VGND VPWR VPWR _14526_/X sky130_fd_sc_hd__o22a_1
X_12787_ _12727_/Y _12785_/X _12786_/Y VGND VGND VPWR VPWR _12787_/X sky130_fd_sc_hd__o21a_1
X_11738_ _10226_/X _11748_/B _10226_/A _11748_/B VGND VGND VPWR VPWR _11746_/A sky130_fd_sc_hd__a2bb2o_1
X_14457_ _13609_/Y _13615_/A _13616_/Y VGND VGND VPWR VPWR _14457_/Y sky130_fd_sc_hd__o21ai_1
X_11669_ _09199_/Y _11666_/Y _09199_/A _11666_/A _11668_/X VGND VGND VPWR VPWR _13132_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14388_ _14329_/X _14386_/X _15612_/B VGND VGND VPWR VPWR _14388_/X sky130_fd_sc_hd__o21a_1
X_13408_ _15470_/A _13348_/B _13348_/Y VGND VGND VPWR VPWR _13408_/X sky130_fd_sc_hd__a21o_1
X_16127_ _15990_/X _16056_/X _15992_/B VGND VGND VPWR VPWR _16127_/X sky130_fd_sc_hd__o21a_1
X_13339_ _13278_/A _13338_/Y _13278_/A _13338_/Y VGND VGND VPWR VPWR _13340_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16058_ _16125_/A _16125_/B VGND VGND VPWR VPWR _16058_/X sky130_fd_sc_hd__and2_1
XFILLER_130_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15009_ _12090_/X _15005_/X _12090_/X _15005_/X VGND VGND VPWR VPWR _15044_/B sky130_fd_sc_hd__a2bb2o_1
X_08880_ _08982_/A _08982_/B VGND VGND VPWR VPWR _08880_/X sky130_fd_sc_hd__and2_1
XFILLER_96_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09501_ _08839_/A _09461_/X _08839_/A _09461_/X VGND VGND VPWR VPWR _09502_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09432_ _09432_/A _09432_/B VGND VGND VPWR VPWR _09432_/X sky130_fd_sc_hd__or2_1
XFILLER_80_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09363_ _08753_/Y _09337_/Y _08753_/Y _09337_/Y VGND VGND VPWR VPWR _11577_/A sky130_fd_sc_hd__a2bb2o_2
X_08314_ _08314_/A VGND VGND VPWR VPWR _08314_/Y sky130_fd_sc_hd__inv_2
X_09294_ _09502_/A _09006_/Y _09540_/A _09231_/Y VGND VGND VPWR VPWR _09294_/X sky130_fd_sc_hd__a31o_1
X_08245_ input5/X _08245_/B VGND VGND VPWR VPWR _08312_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10971_ _11607_/A _10971_/B VGND VGND VPWR VPWR _10972_/A sky130_fd_sc_hd__or2_1
XFILLER_16_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13690_ _14492_/A _13690_/B VGND VGND VPWR VPWR _13690_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12710_ _12707_/A _12707_/B _12707_/Y _12709_/X VGND VGND VPWR VPWR _12710_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12641_ _14170_/A _12639_/X _12640_/X VGND VGND VPWR VPWR _12642_/A sky130_fd_sc_hd__o21ai_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12572_ _14912_/A _12341_/B _12341_/Y VGND VGND VPWR VPWR _12573_/A sky130_fd_sc_hd__o21ai_1
X_15360_ _15296_/X _15360_/B VGND VGND VPWR VPWR _15360_/Y sky130_fd_sc_hd__nand2b_1
X_14311_ _15964_/A _14393_/B VGND VGND VPWR VPWR _14311_/X sky130_fd_sc_hd__and2_1
X_15291_ _15234_/A _15234_/B _15234_/Y VGND VGND VPWR VPWR _15291_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11523_ _10037_/X _11523_/B VGND VGND VPWR VPWR _11523_/X sky130_fd_sc_hd__and2b_1
X_14242_ _14242_/A _14242_/B VGND VGND VPWR VPWR _14371_/B sky130_fd_sc_hd__nor2_1
X_11454_ _12351_/A VGND VGND VPWR VPWR _15540_/A sky130_fd_sc_hd__buf_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10405_ _10405_/A VGND VGND VPWR VPWR _11783_/A sky130_fd_sc_hd__buf_1
XFILLER_125_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14173_ _13443_/A _14132_/A _14130_/Y VGND VGND VPWR VPWR _14173_/Y sky130_fd_sc_hd__a21oi_1
X_11385_ _11259_/X _11384_/Y _11259_/X _11384_/Y VGND VGND VPWR VPWR _11386_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13124_ _13047_/Y _13122_/X _13123_/Y VGND VGND VPWR VPWR _13124_/X sky130_fd_sc_hd__o21a_1
X_10336_ _11727_/A _10335_/B _10335_/Y VGND VGND VPWR VPWR _10336_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13055_ _13055_/A _13029_/X VGND VGND VPWR VPWR _13055_/X sky130_fd_sc_hd__or2b_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _10288_/B VGND VGND VPWR VPWR _10268_/A sky130_fd_sc_hd__inv_2
X_12006_ _11986_/X _12005_/X _11986_/X _12005_/X VGND VGND VPWR VPWR _12073_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10198_ _10197_/Y _10134_/X _10197_/Y _10134_/X VGND VGND VPWR VPWR _10198_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13957_ _15416_/A _13957_/B VGND VGND VPWR VPWR _13957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12908_ _14460_/A _12928_/B VGND VGND VPWR VPWR _12908_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15627_ _16036_/A VGND VGND VPWR VPWR _15673_/A sky130_fd_sc_hd__inv_2
X_13888_ _15420_/A _13961_/B VGND VGND VPWR VPWR _13888_/Y sky130_fd_sc_hd__nor2_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12839_ _15084_/A _12839_/B VGND VGND VPWR VPWR _12839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _15555_/X _15557_/Y _15555_/X _15557_/Y VGND VGND VPWR VPWR _15558_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15489_ _15437_/A _15437_/B _15437_/A _15437_/B VGND VGND VPWR VPWR _15489_/X sky130_fd_sc_hd__a2bb2o_1
X_14509_ _15211_/A _14509_/B VGND VGND VPWR VPWR _14509_/X sky130_fd_sc_hd__or2_1
Xinput30 wbs_dat_i[6] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__buf_1
XFILLER_128_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09981_ _09981_/A _09981_/B VGND VGND VPWR VPWR _09981_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08932_ _10228_/B _08932_/B VGND VGND VPWR VPWR _08932_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08863_ _08795_/X _08801_/A _08803_/Y _08862_/X VGND VGND VPWR VPWR _08863_/X sky130_fd_sc_hd__o22a_1
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08794_ _08794_/A VGND VGND VPWR VPWR _09492_/A sky130_fd_sc_hd__buf_1
XFILLER_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09415_ _09415_/A _09415_/B VGND VGND VPWR VPWR _09415_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09346_ _09346_/A VGND VGND VPWR VPWR _09346_/Y sky130_fd_sc_hd__inv_2
X_09277_ _09256_/X _08910_/Y _09256_/X _08910_/Y VGND VGND VPWR VPWR _10254_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11170_ _12195_/A _11170_/B VGND VGND VPWR VPWR _11170_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10121_ _10120_/X _08989_/Y _10120_/X _08989_/Y VGND VGND VPWR VPWR _10237_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10052_ _10052_/A _10077_/B VGND VGND VPWR VPWR _10052_/X sky130_fd_sc_hd__and2_1
XFILLER_130_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14860_ _14829_/X _14859_/X _14829_/X _14859_/X VGND VGND VPWR VPWR _14930_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14791_ _15455_/A VGND VGND VPWR VPWR _14794_/A sky130_fd_sc_hd__buf_1
X_13811_ _14614_/A _13851_/B VGND VGND VPWR VPWR _13811_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13742_ _13689_/X _13741_/Y _13689_/X _13741_/Y VGND VGND VPWR VPWR _13760_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10954_ _10953_/A _10953_/B _10953_/X _10799_/X VGND VGND VPWR VPWR _10954_/X sky130_fd_sc_hd__o22a_1
XFILLER_16_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16461_ _16357_/A _16461_/D VGND VGND VPWR VPWR _16461_/Q sky130_fd_sc_hd__dfxtp_1
X_10885_ _10774_/X _10884_/Y _10774_/X _10884_/Y VGND VGND VPWR VPWR _10886_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13673_ _15140_/A _13605_/B _13605_/Y VGND VGND VPWR VPWR _13673_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16392_ _16392_/A _16392_/B _16392_/C VGND VGND VPWR VPWR _16454_/A sky130_fd_sc_hd__or3_1
X_12624_ _12624_/A _12624_/B VGND VGND VPWR VPWR _12624_/X sky130_fd_sc_hd__or2_1
X_15412_ _15412_/A _15412_/B VGND VGND VPWR VPWR _15412_/X sky130_fd_sc_hd__or2_1
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12555_ _12628_/A _12628_/B VGND VGND VPWR VPWR _14201_/A sky130_fd_sc_hd__and2_1
X_15343_ _15343_/A _15343_/B VGND VGND VPWR VPWR _15343_/X sky130_fd_sc_hd__or2_1
XFILLER_8_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11506_ _11506_/A _11506_/B VGND VGND VPWR VPWR _11506_/X sky130_fd_sc_hd__and2_1
X_12486_ _13132_/A _12488_/B VGND VGND VPWR VPWR _12486_/Y sky130_fd_sc_hd__nor2_1
X_15274_ _14575_/A _15264_/B _15264_/Y _15273_/Y VGND VGND VPWR VPWR _15274_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14225_ _12594_/X _14225_/B VGND VGND VPWR VPWR _14225_/Y sky130_fd_sc_hd__nand2b_1
X_11437_ _15524_/A _11437_/B VGND VGND VPWR VPWR _11437_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14156_ _14244_/A VGND VGND VPWR VPWR _14230_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11368_ _11572_/A _11368_/B VGND VGND VPWR VPWR _12308_/A sky130_fd_sc_hd__or2_1
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13107_ _15261_/A _13107_/B VGND VGND VPWR VPWR _13107_/Y sky130_fd_sc_hd__nand2_1
X_10319_ _13524_/A _10319_/B VGND VGND VPWR VPWR _10319_/X sky130_fd_sc_hd__and2_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14090_/A _14090_/B VGND VGND VPWR VPWR _14087_/X sky130_fd_sc_hd__and2_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11299_ _11299_/A VGND VGND VPWR VPWR _11299_/Y sky130_fd_sc_hd__inv_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _14976_/A _13127_/B VGND VGND VPWR VPWR _13038_/Y sky130_fd_sc_hd__nor2_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14989_ _14956_/A _14956_/B _14956_/Y _14959_/X VGND VGND VPWR VPWR _14989_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_35_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09200_ _09196_/Y _09199_/A _09198_/X _09199_/Y VGND VGND VPWR VPWR _09200_/X sky130_fd_sc_hd__a22o_1
X_09131_ _09424_/A _09131_/B VGND VGND VPWR VPWR _09131_/Y sky130_fd_sc_hd__nand2_1
X_09062_ _08831_/X _09043_/Y _08831_/X _09043_/Y VGND VGND VPWR VPWR _10018_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09964_ _09997_/A _09997_/B VGND VGND VPWR VPWR _09964_/X sky130_fd_sc_hd__and2_1
XFILLER_103_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _09883_/A _09883_/B _09884_/B VGND VGND VPWR VPWR _09903_/A sky130_fd_sc_hd__a21bo_1
X_08915_ _09401_/A VGND VGND VPWR VPWR _09817_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _09826_/B VGND VGND VPWR VPWR _08847_/A sky130_fd_sc_hd__inv_2
XFILLER_57_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08777_ _10011_/A VGND VGND VPWR VPWR _08778_/A sky130_fd_sc_hd__buf_1
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10670_ _10670_/A VGND VGND VPWR VPWR _10670_/Y sky130_fd_sc_hd__inv_2
X_09329_ _09329_/A _09329_/B VGND VGND VPWR VPWR _09329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12340_ _12242_/X _12339_/Y _12242_/X _12339_/Y VGND VGND VPWR VPWR _12571_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12271_ _11145_/A _12178_/A _11316_/B _12270_/Y VGND VGND VPWR VPWR _12272_/A sky130_fd_sc_hd__o22a_1
XFILLER_134_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11222_ _14028_/A VGND VGND VPWR VPWR _14031_/A sky130_fd_sc_hd__buf_1
X_14010_ _13956_/X _14009_/Y _13956_/X _14009_/Y VGND VGND VPWR VPWR _14061_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11153_ _11141_/X _11152_/Y _11141_/X _11152_/Y VGND VGND VPWR VPWR _11314_/A sky130_fd_sc_hd__o2bb2a_1
X_15961_ _15927_/X _15959_/X _16005_/B VGND VGND VPWR VPWR _15961_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11084_ _13917_/A _11084_/B VGND VGND VPWR VPWR _11084_/X sky130_fd_sc_hd__or2_1
XFILLER_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10104_ _10103_/A _10103_/B _10123_/B VGND VGND VPWR VPWR _10177_/A sky130_fd_sc_hd__o21ai_2
X_15892_ _15892_/A _15892_/B VGND VGND VPWR VPWR _15892_/Y sky130_fd_sc_hd__nand2_1
X_14912_ _14912_/A _14912_/B VGND VGND VPWR VPWR _14912_/Y sky130_fd_sc_hd__nand2_1
X_10035_ _10035_/A _10035_/B VGND VGND VPWR VPWR _10035_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14843_ _14838_/X _14842_/X _14838_/X _14842_/X VGND VGND VPWR VPWR _14944_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14774_ _14774_/A _14774_/B VGND VGND VPWR VPWR _14774_/X sky130_fd_sc_hd__and2_1
XFILLER_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11986_ _13547_/A _11985_/B _11985_/X _11915_/X VGND VGND VPWR VPWR _11986_/X sky130_fd_sc_hd__o22a_1
XFILLER_90_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13725_ _13772_/A _13772_/B VGND VGND VPWR VPWR _13803_/A sky130_fd_sc_hd__and2_1
X_10937_ _13053_/A VGND VGND VPWR VPWR _12103_/A sky130_fd_sc_hd__buf_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16444_ _16434_/A _16434_/B _16434_/Y _16439_/X _16443_/Y VGND VGND VPWR VPWR _16444_/Y
+ sky130_fd_sc_hd__a2111oi_2
X_13656_ _13639_/A _13655_/Y _13639_/A _13655_/Y VGND VGND VPWR VPWR _13700_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12607_ _11422_/X _12607_/B VGND VGND VPWR VPWR _12608_/B sky130_fd_sc_hd__and2b_1
X_10868_ _11974_/A _10724_/B _10724_/Y VGND VGND VPWR VPWR _10868_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16375_ _16320_/A _16320_/B _16320_/Y VGND VGND VPWR VPWR _16375_/Y sky130_fd_sc_hd__o21ai_1
X_13587_ _13547_/A _13547_/B _13548_/A VGND VGND VPWR VPWR _13587_/Y sky130_fd_sc_hd__o21ai_1
X_10799_ _10666_/X _10798_/B _10798_/X _10662_/X VGND VGND VPWR VPWR _10799_/X sky130_fd_sc_hd__o22a_1
XFILLER_129_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12538_ _14113_/A VGND VGND VPWR VPWR _13437_/A sky130_fd_sc_hd__buf_1
X_15326_ _15331_/A _15331_/B VGND VGND VPWR VPWR _15326_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12469_ _12466_/X _12467_/X _12476_/B VGND VGND VPWR VPWR _12469_/X sky130_fd_sc_hd__o21a_1
X_15257_ _15220_/X _15256_/Y _15220_/X _15256_/Y VGND VGND VPWR VPWR _15258_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14208_ _12625_/X _14207_/X _12625_/X _14207_/X VGND VGND VPWR VPWR _14262_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15188_ _15122_/A _15122_/B _15122_/Y VGND VGND VPWR VPWR _15188_/Y sky130_fd_sc_hd__o21ai_1
X_14139_ _14133_/X _14136_/Y _14864_/A _14138_/Y VGND VGND VPWR VPWR _14139_/X sky130_fd_sc_hd__o22a_1
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ _08239_/Y _08699_/A _08239_/A _08699_/Y VGND VGND VPWR VPWR _08701_/B sky130_fd_sc_hd__o22a_1
X_09680_ _09680_/A _09829_/B VGND VGND VPWR VPWR _09683_/A sky130_fd_sc_hd__or2_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08631_ _09225_/B VGND VGND VPWR VPWR _08631_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08562_ _08561_/A _08333_/Y _08561_/Y _08333_/A VGND VGND VPWR VPWR _08563_/B sky130_fd_sc_hd__o22a_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08493_ _08316_/A _08248_/B _08471_/Y _08527_/A VGND VGND VPWR VPWR _08516_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09114_ _09110_/Y _09112_/Y _09113_/Y VGND VGND VPWR VPWR _09118_/B sky130_fd_sc_hd__o21ai_1
X_09045_ _08716_/A _08716_/B _08716_/X _09044_/X VGND VGND VPWR VPWR _09045_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09947_ _09947_/A VGND VGND VPWR VPWR _09947_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09868_/X _08781_/Y _09868_/X _08781_/Y VGND VGND VPWR VPWR _09885_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08829_ _09225_/A _09457_/B _08717_/X VGND VGND VPWR VPWR _08830_/A sky130_fd_sc_hd__o21ai_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11840_ _11840_/A _11840_/B VGND VGND VPWR VPWR _11840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11771_ _12770_/A _11802_/A _11770_/Y VGND VGND VPWR VPWR _11771_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10722_ _13694_/A _10645_/B _10645_/Y VGND VGND VPWR VPWR _10722_/Y sky130_fd_sc_hd__o21ai_1
X_13510_ _13512_/A VGND VGND VPWR VPWR _15040_/A sky130_fd_sc_hd__buf_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14463_/X _14489_/Y _14463_/X _14489_/Y VGND VGND VPWR VPWR _14515_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13441_ _13441_/A _13441_/B VGND VGND VPWR VPWR _13441_/Y sky130_fd_sc_hd__nand2_1
X_10653_ _11980_/A VGND VGND VPWR VPWR _13698_/A sky130_fd_sc_hd__buf_1
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16160_ _16160_/A _16160_/B VGND VGND VPWR VPWR _16268_/B sky130_fd_sc_hd__or2_1
X_13372_ _13313_/A _13313_/B _13313_/X _13371_/X VGND VGND VPWR VPWR _13372_/X sky130_fd_sc_hd__o22a_1
X_10584_ _11910_/A _10648_/B VGND VGND VPWR VPWR _10584_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16091_ _16091_/A _16094_/B VGND VGND VPWR VPWR _16091_/Y sky130_fd_sc_hd__nor2_1
X_12323_ _14081_/A _12320_/B _12321_/Y _12610_/A VGND VGND VPWR VPWR _12324_/B sky130_fd_sc_hd__o22a_1
X_15111_ _15054_/A _15054_/B _15054_/Y VGND VGND VPWR VPWR _15111_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15042_ _15042_/A _15042_/B VGND VGND VPWR VPWR _15042_/X sky130_fd_sc_hd__or2_1
X_12254_ _13048_/A _12254_/B VGND VGND VPWR VPWR _12254_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11205_ _11089_/X _11204_/X _11089_/X _11204_/X VGND VGND VPWR VPWR _11206_/B sky130_fd_sc_hd__a2bb2o_1
X_12185_ _12782_/A _12264_/A _12184_/Y VGND VGND VPWR VPWR _12185_/Y sky130_fd_sc_hd__a21oi_1
X_11136_ _11138_/A VGND VGND VPWR VPWR _11136_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15944_ _15885_/X _15943_/Y _15885_/X _15943_/Y VGND VGND VPWR VPWR _15948_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11067_ _11067_/A _11067_/B VGND VGND VPWR VPWR _11246_/A sky130_fd_sc_hd__or2_1
X_15875_ _15875_/A VGND VGND VPWR VPWR _15890_/A sky130_fd_sc_hd__inv_2
XFILLER_64_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10018_ _10018_/A _10018_/B VGND VGND VPWR VPWR _10061_/B sky130_fd_sc_hd__nor2_1
X_14826_ _14778_/A _14778_/B _14778_/X _14825_/X VGND VGND VPWR VPWR _14826_/X sky130_fd_sc_hd__o22a_1
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14757_ _14757_/A _14757_/B VGND VGND VPWR VPWR _14757_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11969_ _11957_/Y _11967_/X _11968_/Y VGND VGND VPWR VPWR _11969_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13708_ _13708_/A VGND VGND VPWR VPWR _13708_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14688_ _14662_/X _14687_/Y _14662_/X _14687_/Y VGND VGND VPWR VPWR _14740_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16427_ _16412_/Y _16415_/X _16416_/Y _16420_/X _16426_/X VGND VGND VPWR VPWR _16445_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13639_ _13639_/A VGND VGND VPWR VPWR _13639_/Y sky130_fd_sc_hd__inv_2
X_16358_ _16358_/A VGND VGND VPWR VPWR _16358_/X sky130_fd_sc_hd__buf_1
XFILLER_9_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15309_ _14583_/A _15252_/B _15252_/Y VGND VGND VPWR VPWR _15309_/Y sky130_fd_sc_hd__o21ai_1
X_16289_ _16265_/X _16288_/Y _16265_/X _16288_/Y VGND VGND VPWR VPWR _16332_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09801_ _09801_/A _09801_/B VGND VGND VPWR VPWR _09844_/A sky130_fd_sc_hd__or2_1
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09732_ _08567_/X _09734_/B _08567_/X _09734_/B VGND VGND VPWR VPWR _09733_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09663_ _09585_/Y _09661_/X _09662_/Y VGND VGND VPWR VPWR _09663_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08614_ _08650_/A _08614_/B VGND VGND VPWR VPWR _09457_/B sky130_fd_sc_hd__or2_1
X_09594_ _09986_/A VGND VGND VPWR VPWR _09987_/A sky130_fd_sc_hd__buf_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08545_ _09740_/A _08567_/B VGND VGND VPWR VPWR _08546_/A sky130_fd_sc_hd__or2_1
X_08476_ input30/X input14/X VGND VGND VPWR VPWR _08476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09028_ _09028_/A VGND VGND VPWR VPWR _09540_/B sky130_fd_sc_hd__inv_2
XFILLER_123_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13990_ _14832_/A _13990_/B VGND VGND VPWR VPWR _13990_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12941_ _12884_/Y _12939_/X _12940_/Y VGND VGND VPWR VPWR _12941_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15660_ _16027_/A VGND VGND VPWR VPWR _15665_/A sky130_fd_sc_hd__inv_2
XFILLER_73_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12872_ _14757_/A _12946_/B VGND VGND VPWR VPWR _12872_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14611_ _14587_/A _14587_/B _14587_/Y VGND VGND VPWR VPWR _14611_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11823_ _11799_/X _11822_/X _11799_/X _11822_/X VGND VGND VPWR VPWR _11844_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15591_ _14392_/X _15590_/Y _14392_/X _15590_/Y VGND VGND VPWR VPWR _15683_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14585_/A _14585_/B VGND VGND VPWR VPWR _14542_/Y sky130_fd_sc_hd__nor2_1
X_11754_ _11752_/X _11754_/B VGND VGND VPWR VPWR _11754_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_14_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11683_/Y _11684_/Y _11683_/Y _11684_/Y VGND VGND VPWR VPWR _11685_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_81_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14473_ _14473_/A _14473_/B VGND VGND VPWR VPWR _14473_/Y sky130_fd_sc_hd__nor2_1
X_10705_ _11980_/A _10784_/B VGND VGND VPWR VPWR _10705_/Y sky130_fd_sc_hd__nand2_1
X_16212_ _16094_/A _16094_/B _16094_/Y VGND VGND VPWR VPWR _16214_/A sky130_fd_sc_hd__o21ai_1
X_13424_ _13358_/X _13423_/X _13358_/X _13423_/X VGND VGND VPWR VPWR _13424_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10636_ _10608_/Y _10633_/Y _10635_/Y VGND VGND VPWR VPWR _10637_/A sky130_fd_sc_hd__o21ai_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16143_ _15820_/X _16142_/X _15820_/X _16142_/X VGND VGND VPWR VPWR _16144_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13355_ _13349_/Y _13402_/A _13354_/X VGND VGND VPWR VPWR _13355_/Y sky130_fd_sc_hd__o21ai_1
X_10567_ _11923_/A _10677_/B _10566_/Y VGND VGND VPWR VPWR _10568_/A sky130_fd_sc_hd__o21ai_2
X_16074_ _16040_/A _16040_/B _16040_/Y VGND VGND VPWR VPWR _16074_/Y sky130_fd_sc_hd__o21ai_1
X_12306_ _14014_/A _12208_/B _12208_/Y VGND VGND VPWR VPWR _12306_/Y sky130_fd_sc_hd__o21ai_1
X_13286_ _13250_/Y _13284_/Y _13285_/Y VGND VGND VPWR VPWR _13287_/A sky130_fd_sc_hd__o21ai_2
XFILLER_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10498_ _10498_/A VGND VGND VPWR VPWR _10498_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12237_ _12237_/A VGND VGND VPWR VPWR _12237_/X sky130_fd_sc_hd__buf_1
X_15025_ _11728_/Y _14997_/X _11728_/Y _14997_/X VGND VGND VPWR VPWR _15028_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12168_ _13648_/A _12167_/B _12167_/X _12076_/X VGND VGND VPWR VPWR _12168_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12099_ _12074_/X _12098_/Y _12074_/X _12098_/Y VGND VGND VPWR VPWR _12162_/B sky130_fd_sc_hd__a2bb2o_1
X_11119_ _11119_/A VGND VGND VPWR VPWR _11119_/Y sky130_fd_sc_hd__inv_2
X_15927_ _15960_/A _15960_/B VGND VGND VPWR VPWR _15927_/X sky130_fd_sc_hd__and2_1
Xinput6 wbs_adr_i[13] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15858_ _14183_/X _15848_/X _14183_/X _15848_/X VGND VGND VPWR VPWR _15902_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15789_ _15666_/X _15788_/Y _15666_/X _15788_/Y VGND VGND VPWR VPWR _15789_/Y sky130_fd_sc_hd__a2bb2oi_2
X_14809_ _14809_/A _14809_/B VGND VGND VPWR VPWR _14809_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08330_ _08328_/Y _08329_/A _08328_/A _08329_/Y _08304_/A VGND VGND VPWR VPWR _08565_/B
+ sky130_fd_sc_hd__o221a_1
X_08261_ input14/X VGND VGND VPWR VPWR _08341_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_32_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09715_ _09409_/A _09713_/A _10216_/A _09714_/Y VGND VGND VPWR VPWR _09717_/B sky130_fd_sc_hd__o22a_1
XFILLER_67_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09646_ _09642_/Y _10735_/A _09645_/Y VGND VGND VPWR VPWR _09650_/B sky130_fd_sc_hd__o21ai_1
XFILLER_70_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _08692_/A _09154_/A _09528_/A VGND VGND VPWR VPWR _09577_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08527_/A _08318_/Y _08527_/Y _08318_/A VGND VGND VPWR VPWR _08529_/B sky130_fd_sc_hd__o22a_1
XFILLER_23_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08459_ _08459_/A VGND VGND VPWR VPWR _08459_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11470_ _11470_/A VGND VGND VPWR VPWR _11470_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10421_ _10421_/A _10421_/B VGND VGND VPWR VPWR _10422_/A sky130_fd_sc_hd__or2_1
XFILLER_124_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13140_ _15289_/A _13139_/B _13139_/Y VGND VGND VPWR VPWR _13140_/X sky130_fd_sc_hd__a21o_1
X_10352_ _10352_/A _10623_/A VGND VGND VPWR VPWR _10423_/A sky130_fd_sc_hd__nand2_1
X_13071_ _13022_/X _13070_/X _13022_/X _13070_/X VGND VGND VPWR VPWR _13113_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12022_ _11976_/A _11976_/B _11976_/Y VGND VGND VPWR VPWR _12022_/Y sky130_fd_sc_hd__o21ai_1
X_10283_ _10282_/A _11724_/A _10282_/Y _10283_/B2 VGND VGND VPWR VPWR _13478_/B sky130_fd_sc_hd__o22a_1
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13973_ _13972_/A _13972_/B _13972_/Y VGND VGND VPWR VPWR _13973_/X sky130_fd_sc_hd__a21o_1
X_15712_ _16123_/A _15821_/B VGND VGND VPWR VPWR _15712_/X sky130_fd_sc_hd__and2_1
X_12924_ _12924_/A VGND VGND VPWR VPWR _12924_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15643_ _16032_/A VGND VGND VPWR VPWR _15669_/A sky130_fd_sc_hd__inv_2
XFILLER_92_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12855_ _12855_/A _12855_/B VGND VGND VPWR VPWR _12855_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15574_ _15551_/X _15573_/X _15551_/X _15573_/X VGND VGND VPWR VPWR _15575_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12786_/A _12786_/B VGND VGND VPWR VPWR _12786_/Y sky130_fd_sc_hd__nand2_1
X_11806_ _11806_/A _11806_/B VGND VGND VPWR VPWR _11806_/X sky130_fd_sc_hd__or2_1
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14473_/A _14473_/B _14470_/X _14473_/Y VGND VGND VPWR VPWR _14525_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11737_ _11736_/A _11736_/B _10213_/B _11736_/X VGND VGND VPWR VPWR _11748_/B sky130_fd_sc_hd__a22o_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14456_ _14458_/A _14458_/B VGND VGND VPWR VPWR _14456_/Y sky130_fd_sc_hd__nor2_1
X_11668_ _11667_/A _11667_/B _09189_/A _09190_/B _11667_/Y VGND VGND VPWR VPWR _11668_/X
+ sky130_fd_sc_hd__o32a_1
X_14387_ _14387_/A _15958_/A VGND VGND VPWR VPWR _15612_/B sky130_fd_sc_hd__or2_1
X_13407_ _14901_/A _13407_/B VGND VGND VPWR VPWR _13407_/X sky130_fd_sc_hd__and2_1
X_10619_ _13609_/A _10523_/B _10523_/Y VGND VGND VPWR VPWR _10619_/Y sky130_fd_sc_hd__a21oi_1
X_11599_ _11599_/A1 _11598_/Y _11599_/B1 _11598_/A _10959_/X VGND VGND VPWR VPWR _15163_/A
+ sky130_fd_sc_hd__o221a_2
X_16126_ _16058_/X _16124_/X _16386_/B VGND VGND VPWR VPWR _16126_/Y sky130_fd_sc_hd__o21ai_1
X_13338_ _14726_/A _13279_/B _13279_/Y VGND VGND VPWR VPWR _13338_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16057_ _15992_/Y _16056_/X _15992_/Y _16056_/X VGND VGND VPWR VPWR _16125_/B sky130_fd_sc_hd__a2bb2o_1
X_13269_ _15087_/A VGND VGND VPWR VPWR _14721_/A sky130_fd_sc_hd__buf_1
X_15008_ _15046_/A _15046_/B VGND VGND VPWR VPWR _15055_/A sky130_fd_sc_hd__and2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09500_ _09500_/A _09500_/B VGND VGND VPWR VPWR _09500_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09431_ _09431_/A _09431_/B VGND VGND VPWR VPWR _09431_/X sky130_fd_sc_hd__or2_1
XFILLER_52_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09362_ _09362_/A VGND VGND VPWR VPWR _09429_/B sky130_fd_sc_hd__inv_2
X_08313_ _08313_/A VGND VGND VPWR VPWR _08313_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09293_ _09292_/A _09292_/B _08929_/A _09292_/Y VGND VGND VPWR VPWR _09297_/B sky130_fd_sc_hd__o2bb2a_1
X_08244_ input21/X VGND VGND VPWR VPWR _08245_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10970_ _10080_/X _10969_/X _10080_/X _10969_/X VGND VGND VPWR VPWR _10971_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09629_ _09629_/A _09629_/B _09707_/A VGND VGND VPWR VPWR _09629_/X sky130_fd_sc_hd__and3_1
X_12640_ _12640_/A _12640_/B VGND VGND VPWR VPWR _12640_/X sky130_fd_sc_hd__or2_1
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14310_ _14273_/A _14309_/Y _14273_/A _14309_/Y VGND VGND VPWR VPWR _14393_/B sky130_fd_sc_hd__a2bb2o_1
X_12571_ _12571_/A VGND VGND VPWR VPWR _12571_/Y sky130_fd_sc_hd__inv_2
X_15290_ _15289_/A _15289_/B _15289_/Y VGND VGND VPWR VPWR _15290_/X sky130_fd_sc_hd__a21o_1
X_11522_ _11521_/Y _11317_/X _11326_/Y VGND VGND VPWR VPWR _11522_/X sky130_fd_sc_hd__o21a_1
X_14241_ _14242_/A _14242_/B VGND VGND VPWR VPWR _14371_/A sky130_fd_sc_hd__and2_1
XFILLER_109_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11453_ _11258_/X _11452_/Y _11258_/X _11452_/Y VGND VGND VPWR VPWR _12546_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14172_ _15910_/A _14287_/B VGND VGND VPWR VPWR _14172_/X sky130_fd_sc_hd__and2_1
X_10404_ _10402_/A _10403_/A _10402_/Y _10403_/Y _09391_/A VGND VGND VPWR VPWR _10405_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11384_ _14055_/A _11206_/B _11206_/Y VGND VGND VPWR VPWR _11384_/Y sky130_fd_sc_hd__o21ai_1
X_13123_ _15237_/A _13123_/B VGND VGND VPWR VPWR _13123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10335_ _11727_/A _10335_/B VGND VGND VPWR VPWR _10335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13054_ _13772_/A VGND VGND VPWR VPWR _15243_/A sky130_fd_sc_hd__buf_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _09343_/X _10265_/X _09343_/X _10265_/X VGND VGND VPWR VPWR _10288_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12005_ _11009_/A _12075_/B _11009_/A _12075_/B VGND VGND VPWR VPWR _12005_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10197_ _10120_/X _08989_/Y _08468_/Y VGND VGND VPWR VPWR _10197_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_19_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13956_ _13900_/Y _13954_/X _13955_/Y VGND VGND VPWR VPWR _13956_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13887_ _13860_/X _13886_/Y _13860_/X _13886_/Y VGND VGND VPWR VPWR _13961_/B sky130_fd_sc_hd__a2bb2o_1
X_12907_ _12840_/X _12906_/Y _12840_/X _12906_/Y VGND VGND VPWR VPWR _12928_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ _15624_/A _15625_/A _15624_/Y _15625_/Y _15571_/A VGND VGND VPWR VPWR _16036_/A
+ sky130_fd_sc_hd__a221o_2
X_12838_ _15087_/A _12837_/B _12836_/X _12837_/X VGND VGND VPWR VPWR _12838_/X sky130_fd_sc_hd__o22a_1
XFILLER_62_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15556_/Y _15229_/Y _15174_/Y VGND VGND VPWR VPWR _15557_/Y sky130_fd_sc_hd__o21ai_1
X_12769_ _12754_/Y _12767_/X _12768_/Y VGND VGND VPWR VPWR _12769_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15488_ _15554_/A _15554_/B VGND VGND VPWR VPWR _15488_/Y sky130_fd_sc_hd__nor2_1
X_14508_ _15216_/A _14507_/B _13009_/Y _14507_/Y VGND VGND VPWR VPWR _14508_/X sky130_fd_sc_hd__o2bb2a_1
Xinput20 wbs_dat_i[11] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_4
X_14439_ _14438_/A _14438_/B _14438_/Y VGND VGND VPWR VPWR _14439_/X sky130_fd_sc_hd__a21o_1
Xinput31 wbs_dat_i[7] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16109_ _16076_/X _16107_/X _16179_/B VGND VGND VPWR VPWR _16109_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09980_ _09980_/A _09981_/B VGND VGND VPWR VPWR _09980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08931_ _08931_/A VGND VGND VPWR VPWR _08931_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08862_ _09494_/A _08809_/Y _08810_/Y _08861_/X VGND VGND VPWR VPWR _08862_/X sky130_fd_sc_hd__o22a_1
XFILLER_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08793_ _10013_/A _08793_/B VGND VGND VPWR VPWR _08793_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09414_ _09415_/A _09415_/B VGND VGND VPWR VPWR _09414_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09345_ _09561_/A _09345_/B VGND VGND VPWR VPWR _09346_/A sky130_fd_sc_hd__or2_1
X_09276_ _09240_/X _09275_/X _09240_/X _09275_/X VGND VGND VPWR VPWR _10437_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10120_ _10120_/A _10120_/B VGND VGND VPWR VPWR _10120_/X sky130_fd_sc_hd__or2_1
X_10051_ _10024_/X _10050_/Y _10024_/X _10050_/Y VGND VGND VPWR VPWR _10077_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14790_ _14790_/A _14790_/B VGND VGND VPWR VPWR _14790_/X sky130_fd_sc_hd__and2_1
X_13810_ _13767_/X _13809_/X _13767_/X _13809_/X VGND VGND VPWR VPWR _13851_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13741_ _14492_/A _13690_/B _13690_/Y VGND VGND VPWR VPWR _13741_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10953_ _10953_/A _10953_/B VGND VGND VPWR VPWR _10953_/X sky130_fd_sc_hd__and2_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16460_ _16357_/A _16460_/D VGND VGND VPWR VPWR _16460_/Q sky130_fd_sc_hd__dfxtp_1
X_10884_ _13083_/A _10741_/B _10741_/Y VGND VGND VPWR VPWR _10884_/Y sky130_fd_sc_hd__o21ai_1
X_13672_ _13672_/A _13690_/B VGND VGND VPWR VPWR _13672_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16391_ _16389_/X _16390_/Y _16389_/X _16390_/Y VGND VGND VPWR VPWR _16392_/C sky130_fd_sc_hd__a2bb2o_1
X_12623_ _14219_/A _12621_/X _12622_/X VGND VGND VPWR VPWR _12623_/X sky130_fd_sc_hd__o21a_1
X_15411_ _15450_/A _15409_/X _15410_/X VGND VGND VPWR VPWR _15411_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12554_ _12551_/Y _12553_/Y _12551_/A _12553_/A _12503_/A VGND VGND VPWR VPWR _12628_/B
+ sky130_fd_sc_hd__o221a_1
X_15342_ _15375_/A _15340_/X _15341_/X VGND VGND VPWR VPWR _15342_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15273_ _15324_/A _15271_/X _15272_/X VGND VGND VPWR VPWR _15273_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11505_ _12390_/A VGND VGND VPWR VPWR _13974_/A sky130_fd_sc_hd__clkbuf_2
X_14224_ _14230_/A _14224_/B VGND VGND VPWR VPWR _15878_/A sky130_fd_sc_hd__or2_1
X_12485_ _12479_/Y _12484_/Y _12479_/Y _12484_/Y VGND VGND VPWR VPWR _12488_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11436_ _13397_/A VGND VGND VPWR VPWR _15524_/A sky130_fd_sc_hd__buf_1
X_14155_ _14074_/X _14154_/Y _14074_/X _14154_/Y VGND VGND VPWR VPWR _14244_/A sky130_fd_sc_hd__a2bb2o_4
X_11367_ _08977_/X _11366_/X _08977_/X _11366_/X VGND VGND VPWR VPWR _11368_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_125_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14086_ _14901_/A _14083_/B _14083_/X _14085_/Y VGND VGND VPWR VPWR _14090_/B sky130_fd_sc_hd__o22a_1
X_13106_ _13092_/Y _13104_/X _13105_/Y VGND VGND VPWR VPWR _13106_/X sky130_fd_sc_hd__o21a_1
X_10318_ _10299_/X _10317_/X _10299_/X _10317_/X VGND VGND VPWR VPWR _10319_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13037_ _12954_/X _13036_/X _12954_/X _13036_/X VGND VGND VPWR VPWR _13127_/B sky130_fd_sc_hd__a2bb2o_1
X_11298_ _11297_/Y _11123_/X _11164_/Y VGND VGND VPWR VPWR _11298_/X sky130_fd_sc_hd__o21a_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _10247_/A _10247_/B _10247_/X _10248_/Y VGND VGND VPWR VPWR _10252_/B sky130_fd_sc_hd__o22ai_2
XFILLER_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14988_ _14979_/X _14987_/X _14979_/X _14987_/X VGND VGND VPWR VPWR _14988_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13939_ _15392_/A _13939_/B VGND VGND VPWR VPWR _13939_/X sky130_fd_sc_hd__or2_1
XFILLER_62_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15609_ _15609_/A VGND VGND VPWR VPWR _15609_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09130_ _09130_/A VGND VGND VPWR VPWR _09130_/Y sky130_fd_sc_hd__inv_2
X_09061_ _08823_/X _09044_/X _08823_/X _09044_/X VGND VGND VPWR VPWR _10017_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09963_ _09963_/A VGND VGND VPWR VPWR _09963_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08914_ _09066_/A VGND VGND VPWR VPWR _09401_/A sky130_fd_sc_hd__inv_2
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09884_/A _09884_/B _09885_/B VGND VGND VPWR VPWR _09908_/A sky130_fd_sc_hd__a21bo_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08944_/A _08719_/B _08719_/Y VGND VGND VPWR VPWR _09826_/B sky130_fd_sc_hd__a21oi_2
XFILLER_57_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08776_ _10131_/A VGND VGND VPWR VPWR _08776_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09328_ _09327_/A _09327_/B _09327_/X VGND VGND VPWR VPWR _09329_/B sky130_fd_sc_hd__a21boi_1
XFILLER_21_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09259_ _10014_/A _08801_/A _10050_/A _09258_/X VGND VGND VPWR VPWR _09259_/X sky130_fd_sc_hd__o22a_1
XFILLER_126_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12270_ _12270_/A _12270_/B VGND VGND VPWR VPWR _12270_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11221_ _13337_/A VGND VGND VPWR VPWR _14028_/A sky130_fd_sc_hd__inv_2
X_11152_ _11152_/A VGND VGND VPWR VPWR _11152_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10103_ _10103_/A _10103_/B VGND VGND VPWR VPWR _10123_/B sky130_fd_sc_hd__nand2_1
XFILLER_122_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15960_ _15960_/A _15960_/B VGND VGND VPWR VPWR _16005_/B sky130_fd_sc_hd__or2_1
XFILLER_110_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11083_ _11229_/A _11081_/X _11082_/X VGND VGND VPWR VPWR _11083_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15891_ _15877_/Y _15889_/X _15890_/Y VGND VGND VPWR VPWR _15891_/X sky130_fd_sc_hd__o21a_1
X_14911_ _14895_/Y _14909_/X _14910_/Y VGND VGND VPWR VPWR _14911_/X sky130_fd_sc_hd__o21a_1
XFILLER_103_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10034_ _10034_/A _10034_/B VGND VGND VPWR VPWR _10034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14842_ _14841_/A _14841_/B _14841_/Y VGND VGND VPWR VPWR _14842_/X sky130_fd_sc_hd__a21o_1
X_14773_ _14741_/X _14772_/X _14741_/X _14772_/X VGND VGND VPWR VPWR _14774_/B sky130_fd_sc_hd__a2bb2o_1
X_11985_ _13547_/A _11985_/B VGND VGND VPWR VPWR _11985_/X sky130_fd_sc_hd__and2_1
XFILLER_17_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13724_ _13701_/X _13723_/X _13701_/X _13723_/X VGND VGND VPWR VPWR _13772_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10936_ _11590_/A _10936_/B VGND VGND VPWR VPWR _13053_/A sky130_fd_sc_hd__or2_2
X_16443_ _16441_/Y _16442_/Y _16441_/Y _16442_/Y VGND VGND VPWR VPWR _16443_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10867_ _10870_/A VGND VGND VPWR VPWR _14622_/A sky130_fd_sc_hd__buf_1
X_13655_ _15122_/A _13641_/B _13641_/Y VGND VGND VPWR VPWR _13655_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _12606_/A _12606_/B _13405_/B VGND VGND VPWR VPWR _14243_/A sky130_fd_sc_hd__and3_1
X_16374_ _16357_/X _16461_/Q _16358_/X _16397_/C _16361_/X VGND VGND VPWR VPWR _16461_/D
+ sky130_fd_sc_hd__o221a_2
X_13586_ _13640_/A _13641_/B VGND VGND VPWR VPWR _13586_/Y sky130_fd_sc_hd__nor2_1
X_10798_ _11016_/A _10798_/B VGND VGND VPWR VPWR _10798_/X sky130_fd_sc_hd__and2_1
XFILLER_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12537_ _12632_/A _12632_/B VGND VGND VPWR VPWR _14189_/A sky130_fd_sc_hd__and2_1
X_15325_ _15271_/X _15324_/X _15271_/X _15324_/X VGND VGND VPWR VPWR _15331_/B sky130_fd_sc_hd__a2bb2o_1
X_12468_ _13988_/A _12468_/B VGND VGND VPWR VPWR _12476_/B sky130_fd_sc_hd__or2_1
X_15256_ _15202_/A _15202_/B _15202_/Y VGND VGND VPWR VPWR _15256_/Y sky130_fd_sc_hd__o21ai_1
X_14207_ _14207_/A _12626_/X VGND VGND VPWR VPWR _14207_/X sky130_fd_sc_hd__or2b_1
X_11419_ _11250_/X _11419_/B VGND VGND VPWR VPWR _11419_/X sky130_fd_sc_hd__and2b_1
X_15187_ _15187_/A _15187_/B VGND VGND VPWR VPWR _15187_/Y sky130_fd_sc_hd__nand2_1
X_14138_ _14138_/A VGND VGND VPWR VPWR _14138_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12399_ _12400_/A _12400_/B VGND VGND VPWR VPWR _12399_/X sky130_fd_sc_hd__and2_1
X_14069_ _11695_/Y _14068_/X _11695_/Y _14068_/X VGND VGND VPWR VPWR _14069_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08630_ _09225_/A VGND VGND VPWR VPWR _10017_/A sky130_fd_sc_hd__buf_1
XFILLER_27_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08561_ _08561_/A VGND VGND VPWR VPWR _08561_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08492_ _08321_/A _08251_/B _08472_/Y _08538_/A VGND VGND VPWR VPWR _08527_/A sky130_fd_sc_hd__o22a_1
XFILLER_90_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09113_ _09717_/A _09113_/B VGND VGND VPWR VPWR _09113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09044_ _08717_/A _08717_/B _08717_/X _09043_/Y VGND VGND VPWR VPWR _09044_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09946_ _09946_/A VGND VGND VPWR VPWR _09946_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09869_/X _08773_/Y _09869_/X _08773_/Y VGND VGND VPWR VPWR _09886_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08828_ _09458_/A VGND VGND VPWR VPWR _09500_/A sky130_fd_sc_hd__buf_1
XFILLER_73_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08759_ _09330_/B VGND VGND VPWR VPWR _10133_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11770_ _12770_/A _11802_/A VGND VGND VPWR VPWR _11770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _11907_/A VGND VGND VPWR VPWR _13694_/A sky130_fd_sc_hd__buf_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13389_/Y _13438_/X _13439_/Y VGND VGND VPWR VPWR _13440_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10652_ _09969_/Y _10651_/A _10077_/A _10651_/Y _10943_/A VGND VGND VPWR VPWR _11980_/A
+ sky130_fd_sc_hd__a221o_2
X_13371_ _13378_/A _13369_/X _13370_/X VGND VGND VPWR VPWR _13371_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10583_ _10534_/X _10582_/Y _10534_/X _10582_/Y VGND VGND VPWR VPWR _10648_/B sky130_fd_sc_hd__a2bb2o_1
X_16090_ _16086_/Y _16223_/A _16089_/Y VGND VGND VPWR VPWR _16094_/B sky130_fd_sc_hd__o21ai_1
X_12322_ _12322_/A _13405_/B VGND VGND VPWR VPWR _12610_/A sky130_fd_sc_hd__or2_1
X_15110_ _15110_/A _15110_/B VGND VGND VPWR VPWR _15110_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12253_ _12292_/A VGND VGND VPWR VPWR _13204_/A sky130_fd_sc_hd__buf_1
X_15041_ _15064_/A _15039_/X _15040_/X VGND VGND VPWR VPWR _15041_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11204_ _11204_/A _11090_/X VGND VGND VPWR VPWR _11204_/X sky130_fd_sc_hd__or2b_1
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12184_ _12782_/A _12264_/A VGND VGND VPWR VPWR _12184_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11135_ _12172_/A VGND VGND VPWR VPWR _13503_/A sky130_fd_sc_hd__buf_1
X_15943_ _15886_/A _15886_/B _15886_/Y VGND VGND VPWR VPWR _15943_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11066_ _12043_/B _11066_/B _13096_/A VGND VGND VPWR VPWR _11067_/B sky130_fd_sc_hd__and3_1
XFILLER_76_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10017_ _10017_/A _10017_/B VGND VGND VPWR VPWR _10065_/B sky130_fd_sc_hd__nor2_1
X_15874_ _15892_/A _15892_/B VGND VGND VPWR VPWR _15874_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14825_ _14782_/A _14782_/B _14782_/X _14824_/X VGND VGND VPWR VPWR _14825_/X sky130_fd_sc_hd__o22a_1
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14756_ _14751_/X _14755_/X _14751_/X _14755_/X VGND VGND VPWR VPWR _14757_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11968_ _11968_/A _11968_/B VGND VGND VPWR VPWR _11968_/Y sky130_fd_sc_hd__nand2_1
X_13707_ _13715_/A VGND VGND VPWR VPWR _15116_/A sky130_fd_sc_hd__buf_1
XFILLER_44_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10919_ _14618_/A _10919_/B VGND VGND VPWR VPWR _10919_/X sky130_fd_sc_hd__or2_1
X_14687_ _15349_/A _14742_/B _14686_/Y VGND VGND VPWR VPWR _14687_/Y sky130_fd_sc_hd__o21ai_1
X_11899_ _11885_/Y _11897_/Y _11898_/Y VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__o21ai_1
XFILLER_32_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16426_ _16426_/A _16434_/A VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__or2b_1
X_13638_ _13589_/Y _13635_/Y _13637_/Y VGND VGND VPWR VPWR _13639_/A sky130_fd_sc_hd__o21ai_1
X_16357_ _16357_/A VGND VGND VPWR VPWR _16357_/X sky130_fd_sc_hd__buf_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13569_ _13529_/A _13529_/B _13529_/Y VGND VGND VPWR VPWR _13569_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15308_ _15343_/A _15343_/B VGND VGND VPWR VPWR _15372_/A sky130_fd_sc_hd__and2_1
XFILLER_8_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16288_ _16266_/A _16332_/A _16266_/Y VGND VGND VPWR VPWR _16288_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15239_ _15226_/X _15238_/Y _15226_/X _15238_/Y VGND VGND VPWR VPWR _15240_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09800_ _09800_/A _09834_/A VGND VGND VPWR VPWR _09801_/B sky130_fd_sc_hd__or2_1
XFILLER_113_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09731_ _09731_/A _09731_/B VGND VGND VPWR VPWR _09734_/B sky130_fd_sc_hd__or2_1
XFILLER_39_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09662_ _09993_/A _09662_/B VGND VGND VPWR VPWR _09662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08613_ _08612_/A _08354_/Y _08612_/Y _08354_/A VGND VGND VPWR VPWR _08614_/B sky130_fd_sc_hd__o22a_1
X_09593_ _09512_/X _09592_/X _09512_/X _09592_/X VGND VGND VPWR VPWR _09986_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _09860_/A VGND VGND VPWR VPWR _09740_/A sky130_fd_sc_hd__inv_2
XFILLER_82_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08475_ input15/X input31/X VGND VGND VPWR VPWR _08475_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09027_ _09005_/Y _08657_/Y _09005_/Y _08657_/Y VGND VGND VPWR VPWR _09028_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09929_ _09347_/B _09924_/Y _09863_/B VGND VGND VPWR VPWR _09929_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12940_ _12940_/A _12940_/B VGND VGND VPWR VPWR _12940_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12871_ _12858_/X _12870_/Y _12858_/X _12870_/Y VGND VGND VPWR VPWR _12946_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14610_ _14610_/A VGND VGND VPWR VPWR _15345_/A sky130_fd_sc_hd__buf_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11822_ _09949_/A _11773_/B _09949_/A _11773_/B VGND VGND VPWR VPWR _11822_/X sky130_fd_sc_hd__a2bb2o_1
X_15590_ _14311_/X _15590_/B VGND VGND VPWR VPWR _15590_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14520_/X _14540_/X _14520_/X _14540_/X VGND VGND VPWR VPWR _14585_/B sky130_fd_sc_hd__a2bb2o_1
X_11753_ _11753_/A _11753_/B VGND VGND VPWR VPWR _11754_/B sky130_fd_sc_hd__or2_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11671_/A _15433_/A _11671_/Y _11576_/Y VGND VGND VPWR VPWR _11684_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_81_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10704_ _10655_/X _10703_/Y _10655_/X _10703_/Y VGND VGND VPWR VPWR _10784_/B sky130_fd_sc_hd__a2bb2o_1
X_14472_ _11932_/Y _14471_/X _11932_/Y _14471_/X VGND VGND VPWR VPWR _14473_/B sky130_fd_sc_hd__o2bb2a_1
X_16211_ _16255_/A _16322_/A VGND VGND VPWR VPWR _16211_/Y sky130_fd_sc_hd__nor2_1
X_13423_ _13337_/A _13337_/B _13337_/A _13337_/B VGND VGND VPWR VPWR _13423_/X sky130_fd_sc_hd__a2bb2o_1
X_10635_ _12997_/A _10635_/B VGND VGND VPWR VPWR _10635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16142_ _15712_/X _16142_/B VGND VGND VPWR VPWR _16142_/X sky130_fd_sc_hd__and2b_1
X_13354_ _15473_/A _13354_/B VGND VGND VPWR VPWR _13354_/X sky130_fd_sc_hd__or2_1
XFILLER_10_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12305_ _12305_/A _12305_/B VGND VGND VPWR VPWR _12305_/Y sky130_fd_sc_hd__nand2_1
X_10566_ _11923_/A _10677_/B VGND VGND VPWR VPWR _10566_/Y sky130_fd_sc_hd__nand2_1
X_16073_ _16110_/A _16110_/B VGND VGND VPWR VPWR _16073_/X sky130_fd_sc_hd__and2_1
X_13285_ _14730_/A _13285_/B VGND VGND VPWR VPWR _13285_/Y sky130_fd_sc_hd__nand2_1
X_10497_ _09838_/A _09838_/B _09839_/A VGND VGND VPWR VPWR _10498_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12236_ _12234_/Y _12235_/X _12234_/Y _12235_/X VGND VGND VPWR VPWR _12238_/B sky130_fd_sc_hd__a2bb2o_1
X_15024_ _15030_/A _15030_/B VGND VGND VPWR VPWR _15079_/A sky130_fd_sc_hd__and2_1
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12167_ _13648_/A _12167_/B VGND VGND VPWR VPWR _12167_/X sky130_fd_sc_hd__and2_1
XFILLER_123_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11118_ _09782_/A _09782_/B _09782_/Y VGND VGND VPWR VPWR _11119_/A sky130_fd_sc_hd__o21ai_1
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12098_ _13705_/A _12165_/B _12097_/Y VGND VGND VPWR VPWR _12098_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15926_ _15897_/X _15925_/Y _15897_/X _15925_/Y VGND VGND VPWR VPWR _15960_/B sky130_fd_sc_hd__a2bb2o_1
Xinput7 wbs_adr_i[14] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_4
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11049_ _12841_/A VGND VGND VPWR VPWR _15081_/A sky130_fd_sc_hd__buf_1
XFILLER_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15857_ _15857_/A VGND VGND VPWR VPWR _15902_/A sky130_fd_sc_hd__inv_2
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14808_ _14723_/X _14807_/X _14723_/X _14807_/X VGND VGND VPWR VPWR _14809_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15788_ _15654_/X _15788_/B VGND VGND VPWR VPWR _15788_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_52_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14739_ _14780_/A _14737_/X _14738_/X VGND VGND VPWR VPWR _14739_/X sky130_fd_sc_hd__o21a_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08260_ input15/X _08260_/B VGND VGND VPWR VPWR _08337_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16409_ _16409_/A VGND VGND VPWR VPWR _16409_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_133_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09714_ _09714_/A _09714_/B VGND VGND VPWR VPWR _09714_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09645_ _09960_/A _09645_/B VGND VGND VPWR VPWR _09645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09515_/X _09575_/X _09515_/X _09575_/X VGND VGND VPWR VPWR _09995_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08527_/A VGND VGND VPWR VPWR _08527_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_51_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08458_ _08532_/B _08453_/Y _09330_/A VGND VGND VPWR VPWR _08459_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10420_ _10906_/A _10420_/B VGND VGND VPWR VPWR _12234_/A sky130_fd_sc_hd__nand2_4
X_08389_ _08389_/A VGND VGND VPWR VPWR _08389_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10351_ _10521_/A VGND VGND VPWR VPWR _10623_/A sky130_fd_sc_hd__inv_2
XFILLER_124_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13070_ _13070_/A _13023_/X VGND VGND VPWR VPWR _13070_/X sky130_fd_sc_hd__or2b_1
X_10282_ _10282_/A VGND VGND VPWR VPWR _10282_/Y sky130_fd_sc_hd__inv_2
X_12021_ _12061_/A VGND VGND VPWR VPWR _13194_/A sky130_fd_sc_hd__buf_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13972_ _13972_/A _13972_/B VGND VGND VPWR VPWR _13972_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15711_ _15695_/X _15710_/Y _15695_/X _15710_/Y VGND VGND VPWR VPWR _15821_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12923_ _13005_/A _12922_/B _12921_/X _12922_/Y VGND VGND VPWR VPWR _12924_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15642_ _15640_/A _15641_/A _15640_/Y _15641_/Y _15571_/A VGND VGND VPWR VPWR _16032_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_74_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12854_ _12805_/Y _12852_/X _12853_/Y VGND VGND VPWR VPWR _12854_/X sky130_fd_sc_hd__o21a_1
X_15573_ _15491_/X _15573_/B VGND VGND VPWR VPWR _15573_/X sky130_fd_sc_hd__and2b_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12785_ _12730_/Y _12783_/X _12784_/Y VGND VGND VPWR VPWR _12785_/X sky130_fd_sc_hd__o21a_1
X_11805_ _11850_/A VGND VGND VPWR VPWR _12772_/A sky130_fd_sc_hd__buf_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14476_/A _14476_/B _14469_/X _14476_/Y VGND VGND VPWR VPWR _14524_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11736_ _11736_/A _11736_/B VGND VGND VPWR VPWR _11736_/X sky130_fd_sc_hd__or2_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14455_ _14430_/X _14454_/X _14430_/X _14454_/X VGND VGND VPWR VPWR _14458_/B sky130_fd_sc_hd__a2bb2o_1
X_11667_ _11667_/A _11667_/B VGND VGND VPWR VPWR _11667_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14386_ _14335_/X _14384_/X _15620_/B VGND VGND VPWR VPWR _14386_/X sky130_fd_sc_hd__o21a_1
X_13406_ _14904_/A _13404_/B _13404_/X _14239_/A VGND VGND VPWR VPWR _13407_/B sky130_fd_sc_hd__o22a_1
X_10618_ _11892_/A VGND VGND VPWR VPWR _13004_/A sky130_fd_sc_hd__buf_1
X_11598_ _11598_/A VGND VGND VPWR VPWR _11598_/Y sky130_fd_sc_hd__inv_2
X_16125_ _16125_/A _16125_/B VGND VGND VPWR VPWR _16386_/B sky130_fd_sc_hd__or2_1
X_13337_ _13337_/A _13337_/B VGND VGND VPWR VPWR _13337_/X sky130_fd_sc_hd__and2_1
X_10549_ _10549_/A VGND VGND VPWR VPWR _10549_/Y sky130_fd_sc_hd__inv_2
X_16056_ _15995_/X _16054_/X _16059_/B VGND VGND VPWR VPWR _16056_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13268_ _13274_/A _13274_/B VGND VGND VPWR VPWR _13268_/Y sky130_fd_sc_hd__nor2_1
X_15007_ _12182_/X _15006_/X _12182_/X _15006_/X VGND VGND VPWR VPWR _15046_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12219_ _12146_/X _12218_/X _12146_/X _12218_/X VGND VGND VPWR VPWR _12220_/B sky130_fd_sc_hd__a2bb2o_1
X_13199_ _13156_/Y _13197_/X _13198_/Y VGND VGND VPWR VPWR _13199_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15909_ _15856_/Y _15907_/X _15908_/Y VGND VGND VPWR VPWR _15909_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09430_ _09430_/A _09430_/B VGND VGND VPWR VPWR _09430_/X sky130_fd_sc_hd__or2_1
XFILLER_37_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09361_ _09360_/X _09357_/X _09360_/X _09357_/X VGND VGND VPWR VPWR _09362_/A sky130_fd_sc_hd__a2bb2o_1
X_08312_ _08312_/A _08312_/B VGND VGND VPWR VPWR _08313_/A sky130_fd_sc_hd__or2_1
X_09292_ _09292_/A _09292_/B VGND VGND VPWR VPWR _09292_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08243_ input5/X VGND VGND VPWR VPWR _08311_/A sky130_fd_sc_hd__inv_2
XFILLER_106_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09628_ _09628_/A _09628_/B VGND VGND VPWR VPWR _09628_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09559_ _08692_/A _09154_/A _09528_/Y _09558_/X VGND VGND VPWR VPWR _09559_/X sky130_fd_sc_hd__o22a_1
X_12570_ _12566_/Y _12569_/Y _12566_/A _12569_/A _11709_/A VGND VGND VPWR VPWR _12624_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11521_ _11521_/A _11521_/B VGND VGND VPWR VPWR _11521_/Y sky130_fd_sc_hd__nor2_1
X_14240_ _14239_/A _14238_/Y _14243_/B _14238_/A _14244_/A VGND VGND VPWR VPWR _14242_/B
+ sky130_fd_sc_hd__a221o_1
X_11452_ _14108_/A _11213_/B _11213_/Y VGND VGND VPWR VPWR _11452_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14171_ _12639_/X _14170_/X _12639_/X _14170_/X VGND VGND VPWR VPWR _14287_/B sky130_fd_sc_hd__a2bb2o_1
X_11383_ _12314_/A VGND VGND VPWR VPWR _14113_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10403_ _10403_/A VGND VGND VPWR VPWR _10403_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13122_ _13052_/Y _13120_/X _13121_/Y VGND VGND VPWR VPWR _13122_/X sky130_fd_sc_hd__o21a_1
X_10334_ _13529_/A VGND VGND VPWR VPWR _15028_/A sky130_fd_sc_hd__buf_1
XFILLER_3_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13053_ _13053_/A VGND VGND VPWR VPWR _13772_/A sky130_fd_sc_hd__inv_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _10197_/Y _10264_/Y _10197_/Y _10264_/Y VGND VGND VPWR VPWR _10265_/X sky130_fd_sc_hd__a2bb2o_1
X_12004_ _12077_/B _12003_/Y _12077_/B _12003_/Y VGND VGND VPWR VPWR _12075_/B sky130_fd_sc_hd__o2bb2a_1
X_10196_ _09341_/X _10195_/Y _09341_/X _10195_/Y VGND VGND VPWR VPWR _10196_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13955_ _15414_/A _13955_/B VGND VGND VPWR VPWR _13955_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13886_ _14832_/A _13990_/B _13885_/Y VGND VGND VPWR VPWR _13886_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12906_ _12841_/A _12841_/B _12841_/Y VGND VGND VPWR VPWR _12906_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _15625_/A VGND VGND VPWR VPWR _15625_/Y sky130_fd_sc_hd__inv_2
X_12837_ _12837_/A _12837_/B VGND VGND VPWR VPWR _12837_/X sky130_fd_sc_hd__and2_1
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _15556_/A _15556_/B VGND VGND VPWR VPWR _15556_/Y sky130_fd_sc_hd__nor2_1
X_12768_ _12768_/A _12768_/B VGND VGND VPWR VPWR _12768_/Y sky130_fd_sc_hd__nand2_1
X_15487_ _15434_/Y _15486_/X _15434_/Y _15486_/X VGND VGND VPWR VPWR _15554_/B sky130_fd_sc_hd__a2bb2o_1
X_14507_ _15216_/A _14507_/B VGND VGND VPWR VPWR _14507_/Y sky130_fd_sc_hd__nor2_1
X_11719_ _11719_/A VGND VGND VPWR VPWR _11720_/B sky130_fd_sc_hd__inv_4
X_12699_ _12699_/A _12699_/B VGND VGND VPWR VPWR _12699_/Y sky130_fd_sc_hd__nor2_1
Xinput21 wbs_dat_i[12] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_4
X_14438_ _14438_/A _14438_/B VGND VGND VPWR VPWR _14438_/Y sky130_fd_sc_hd__nor2_1
Xinput10 wbs_adr_i[2] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_4
Xinput32 wbs_dat_i[8] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__buf_4
X_14369_ _14369_/A VGND VGND VPWR VPWR _15662_/B sky130_fd_sc_hd__inv_6
X_16108_ _16108_/A _16108_/B VGND VGND VPWR VPWR _16179_/B sky130_fd_sc_hd__or2_1
XFILLER_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16039_ _16013_/Y _16037_/X _16038_/Y VGND VGND VPWR VPWR _16039_/X sky130_fd_sc_hd__o21a_1
XFILLER_97_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08930_ _08930_/A _10287_/A VGND VGND VPWR VPWR _08931_/A sky130_fd_sc_hd__or2_2
XFILLER_69_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08861_ _09496_/A _08817_/A _08819_/Y _08860_/X VGND VGND VPWR VPWR _08861_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08792_ _08793_/B VGND VGND VPWR VPWR _08792_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09413_ _09285_/Y _10879_/A _09412_/X VGND VGND VPWR VPWR _09415_/B sky130_fd_sc_hd__o21ai_1
XFILLER_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09344_ _08703_/A _09791_/C _09937_/A _08509_/A VGND VGND VPWR VPWR _09344_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09275_ _08610_/A _09803_/A _09220_/A VGND VGND VPWR VPWR _09275_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10050_ _10050_/A _10050_/B VGND VGND VPWR VPWR _10050_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13740_ _13762_/A _13762_/B VGND VGND VPWR VPWR _13818_/A sky130_fd_sc_hd__and2_1
X_10952_ _12097_/A VGND VGND VPWR VPWR _13705_/A sky130_fd_sc_hd__buf_1
XFILLER_56_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15410_ _15410_/A _15410_/B VGND VGND VPWR VPWR _15410_/X sky130_fd_sc_hd__or2_1
X_10883_ _10886_/A VGND VGND VPWR VPWR _14630_/A sky130_fd_sc_hd__buf_1
XFILLER_71_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13671_ _13619_/X _13670_/Y _13619_/X _13670_/Y VGND VGND VPWR VPWR _13690_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16390_ _16276_/X _16339_/X _16278_/B VGND VGND VPWR VPWR _16390_/Y sky130_fd_sc_hd__o21ai_1
X_12622_ _12622_/A _12622_/B VGND VGND VPWR VPWR _12622_/X sky130_fd_sc_hd__or2_1
X_12553_ _12553_/A VGND VGND VPWR VPWR _12553_/Y sky130_fd_sc_hd__inv_2
X_15341_ _15341_/A _15341_/B VGND VGND VPWR VPWR _15341_/X sky130_fd_sc_hd__or2_1
XFILLER_12_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15272_ _15272_/A _15272_/B VGND VGND VPWR VPWR _15272_/X sky130_fd_sc_hd__or2_1
X_11504_ _12948_/A VGND VGND VPWR VPWR _12390_/A sky130_fd_sc_hd__inv_2
XFILLER_12_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14223_ _14089_/Y _14222_/X _14089_/Y _14222_/X VGND VGND VPWR VPWR _14224_/B sky130_fd_sc_hd__a2bb2oi_1
X_12484_ _13994_/A _12480_/B _12480_/Y VGND VGND VPWR VPWR _12484_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11435_ _11255_/X _11434_/Y _11255_/X _11434_/Y VGND VGND VPWR VPWR _12576_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14154_ _14152_/X _14153_/Y _14152_/X _14153_/Y VGND VGND VPWR VPWR _14154_/Y sky130_fd_sc_hd__a2bb2oi_2
X_11366_ _08890_/X _11366_/B VGND VGND VPWR VPWR _11366_/X sky130_fd_sc_hd__and2b_1
XFILLER_113_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14085_ _14048_/X _14084_/X _14048_/X _14084_/X VGND VGND VPWR VPWR _14085_/Y sky130_fd_sc_hd__a2bb2oi_1
X_13105_ _15264_/A _13105_/B VGND VGND VPWR VPWR _13105_/Y sky130_fd_sc_hd__nand2_1
X_11297_ _12189_/A _11297_/B VGND VGND VPWR VPWR _11297_/Y sky130_fd_sc_hd__nor2_1
X_10317_ _10367_/A _12701_/A _10316_/Y VGND VGND VPWR VPWR _10317_/X sky130_fd_sc_hd__a21o_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _13040_/A _13034_/X _13035_/X VGND VGND VPWR VPWR _13036_/X sky130_fd_sc_hd__o21a_1
X_10248_ _10248_/A VGND VGND VPWR VPWR _10248_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_3_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10179_ _10180_/A _10180_/B VGND VGND VPWR VPWR _10179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14987_ _14981_/X _14986_/X _14981_/X _14986_/X VGND VGND VPWR VPWR _14987_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13938_ _15396_/A _13937_/B _13936_/X _13937_/X VGND VGND VPWR VPWR _13938_/X sky130_fd_sc_hd__o22a_1
XFILLER_93_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13869_ _15104_/A _13497_/B _13497_/Y VGND VGND VPWR VPWR _13869_/Y sky130_fd_sc_hd__o21ai_1
X_15608_ _14916_/A _15540_/B _15540_/Y VGND VGND VPWR VPWR _15609_/A sky130_fd_sc_hd__o21ai_1
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15539_ _15539_/A VGND VGND VPWR VPWR _15539_/Y sky130_fd_sc_hd__clkinvlp_2
X_09060_ _08814_/X _09045_/X _08814_/X _09045_/X VGND VGND VPWR VPWR _10016_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09962_ _09962_/A VGND VGND VPWR VPWR _09962_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08913_ _09041_/A _08913_/B VGND VGND VPWR VPWR _09066_/A sky130_fd_sc_hd__or2_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09885_/A _09885_/B _09886_/B VGND VGND VPWR VPWR _09913_/A sky130_fd_sc_hd__a21bo_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08844_/A _10123_/A VGND VGND VPWR VPWR _08844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08775_ _09332_/B VGND VGND VPWR VPWR _10131_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09327_ _09327_/A _09327_/B VGND VGND VPWR VPWR _09327_/X sky130_fd_sc_hd__or2_1
X_09258_ _08904_/X _08809_/Y _10073_/A _09257_/X VGND VGND VPWR VPWR _09258_/X sky130_fd_sc_hd__o22a_1
X_09189_ _09189_/A VGND VGND VPWR VPWR _09190_/B sky130_fd_sc_hd__inv_2
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11220_ _11220_/A _11220_/B VGND VGND VPWR VPWR _13337_/A sky130_fd_sc_hd__or2_1
XFILLER_107_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11151_ _12270_/A _11316_/B _11150_/Y VGND VGND VPWR VPWR _11152_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10102_ _10102_/A _10102_/B VGND VGND VPWR VPWR _10103_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11082_ _13921_/A _11082_/B VGND VGND VPWR VPWR _11082_/X sky130_fd_sc_hd__or2_1
X_15890_ _15890_/A _15890_/B VGND VGND VPWR VPWR _15890_/Y sky130_fd_sc_hd__nand2_1
X_14910_ _14910_/A _14910_/B VGND VGND VPWR VPWR _14910_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10033_ _09338_/X _10008_/X _10030_/Y _10032_/Y VGND VGND VPWR VPWR _10034_/B sky130_fd_sc_hd__a31o_1
XFILLER_76_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14841_ _14841_/A _14841_/B VGND VGND VPWR VPWR _14841_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14772_ _14772_/A _14771_/X VGND VGND VPWR VPWR _14772_/X sky130_fd_sc_hd__or2b_1
XFILLER_84_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11984_ _11983_/Y _11913_/X _11936_/Y VGND VGND VPWR VPWR _11984_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13723_ _13723_/A _13702_/X VGND VGND VPWR VPWR _13723_/X sky130_fd_sc_hd__or2b_1
XFILLER_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10935_ _09659_/X _10934_/X _09659_/X _10934_/X VGND VGND VPWR VPWR _10936_/B sky130_fd_sc_hd__a2bb2oi_1
X_16442_ _16415_/X _16420_/X _16426_/X VGND VGND VPWR VPWR _16442_/Y sky130_fd_sc_hd__a21boi_1
X_10866_ _12059_/A VGND VGND VPWR VPWR _10870_/A sky130_fd_sc_hd__inv_2
X_13654_ _13702_/A _13702_/B VGND VGND VPWR VPWR _13723_/A sky130_fd_sc_hd__and2_1
XFILLER_44_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16373_ _16321_/X _16372_/Y _16321_/X _16372_/Y VGND VGND VPWR VPWR _16397_/C sky130_fd_sc_hd__a2bb2o_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12605_ _12618_/A _12618_/B VGND VGND VPWR VPWR _14231_/A sky130_fd_sc_hd__and2_1
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15324_ _15324_/A _15272_/X VGND VGND VPWR VPWR _15324_/X sky130_fd_sc_hd__or2b_1
X_10797_ _12007_/A VGND VGND VPWR VPWR _13640_/A sky130_fd_sc_hd__buf_1
X_13585_ _13580_/X _13584_/Y _13580_/X _13584_/Y VGND VGND VPWR VPWR _13641_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12536_ _12535_/A _12535_/B _12535_/Y _12503_/X VGND VGND VPWR VPWR _12632_/B sky130_fd_sc_hd__o211a_1
XFILLER_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12467_ _12399_/X _12361_/X _12401_/B VGND VGND VPWR VPWR _12467_/X sky130_fd_sc_hd__o21a_1
X_15255_ _15255_/A _15255_/B VGND VGND VPWR VPWR _15255_/Y sky130_fd_sc_hd__nand2_1
X_14206_ _14206_/A _14206_/B VGND VGND VPWR VPWR _15869_/A sky130_fd_sc_hd__or2_1
XFILLER_99_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15186_ _15155_/X _15185_/Y _15155_/X _15185_/Y VGND VGND VPWR VPWR _15187_/B sky130_fd_sc_hd__a2bb2o_1
X_11418_ _09403_/X _08931_/A _08931_/Y _10514_/Y _08997_/A VGND VGND VPWR VPWR _13404_/A
+ sky130_fd_sc_hd__o221a_4
X_14137_ _14137_/A VGND VGND VPWR VPWR _14864_/A sky130_fd_sc_hd__inv_2
X_12398_ _12363_/Y _12397_/X _12363_/Y _12397_/X VGND VGND VPWR VPWR _12400_/B sky130_fd_sc_hd__o2bb2a_1
X_11349_ _11482_/A _11482_/B _11482_/A _11482_/B VGND VGND VPWR VPWR _11349_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14068_ _14002_/X _14066_/X _14146_/B VGND VGND VPWR VPWR _14068_/X sky130_fd_sc_hd__o21a_1
X_13019_ _14488_/A _13019_/B VGND VGND VPWR VPWR _13019_/X sky130_fd_sc_hd__or2_1
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08560_ _08688_/A _10117_/B VGND VGND VPWR VPWR _08886_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08491_ _08326_/A _08254_/B _08473_/Y _08549_/A VGND VGND VPWR VPWR _08538_/A sky130_fd_sc_hd__o22a_1
XFILLER_90_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09112_ _09112_/A VGND VGND VPWR VPWR _09112_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09043_ _08718_/Y _09042_/X _08724_/X VGND VGND VPWR VPWR _09043_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09945_ _10252_/A _09309_/B _09309_/Y VGND VGND VPWR VPWR _09947_/A sky130_fd_sc_hd__o21ai_1
XFILLER_112_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09876_ _09870_/X _08765_/Y _09870_/X _08765_/Y VGND VGND VPWR VPWR _09887_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _10017_/A _10125_/A VGND VGND VPWR VPWR _08827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08758_ _08757_/A _08745_/A _08757_/Y _08745_/Y VGND VGND VPWR VPWR _09330_/B sky130_fd_sc_hd__o22a_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08689_ _08886_/A _08687_/X _08886_/B VGND VGND VPWR VPWR _08689_/X sky130_fd_sc_hd__o21ba_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10720_ _13073_/A VGND VGND VPWR VPWR _11974_/A sky130_fd_sc_hd__buf_1
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10651_ _10651_/A VGND VGND VPWR VPWR _10651_/Y sky130_fd_sc_hd__inv_2
X_13370_ _13370_/A _13370_/B VGND VGND VPWR VPWR _13370_/X sky130_fd_sc_hd__or2_1
X_10582_ _13632_/A _10654_/B _10581_/Y VGND VGND VPWR VPWR _10582_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12321_ _12321_/A VGND VGND VPWR VPWR _12321_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12252_ _12251_/Y _12158_/X _12198_/Y VGND VGND VPWR VPWR _12252_/X sky130_fd_sc_hd__o21a_1
X_15040_ _15040_/A _15040_/B VGND VGND VPWR VPWR _15040_/X sky130_fd_sc_hd__or2_1
XFILLER_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11203_ _14055_/A VGND VGND VPWR VPWR _15452_/A sky130_fd_sc_hd__buf_1
XFILLER_5_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12183_ _12268_/B _12182_/X _12268_/B _12182_/X VGND VGND VPWR VPWR _12264_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11134_ _10083_/A _11133_/Y _09966_/Y _11133_/A _10959_/X VGND VGND VPWR VPWR _12172_/A
+ sky130_fd_sc_hd__o221a_1
X_15942_ _15950_/A _15950_/B VGND VGND VPWR VPWR _15942_/X sky130_fd_sc_hd__and2_1
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11065_ _13753_/A _11065_/B VGND VGND VPWR VPWR _13096_/A sky130_fd_sc_hd__or2_1
XFILLER_49_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10016_ _10016_/A _10016_/B VGND VGND VPWR VPWR _10069_/B sky130_fd_sc_hd__nor2_1
X_15873_ _14213_/X _15843_/X _14213_/X _15843_/X VGND VGND VPWR VPWR _15892_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14824_ _14786_/A _14786_/B _14786_/X _14823_/X VGND VGND VPWR VPWR _14824_/X sky130_fd_sc_hd__o22a_1
XFILLER_36_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11967_ _12040_/A _11965_/X _11966_/X VGND VGND VPWR VPWR _11967_/X sky130_fd_sc_hd__o21a_1
X_14755_ _14754_/A _14754_/B _14754_/Y VGND VGND VPWR VPWR _14755_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10918_ _10918_/A VGND VGND VPWR VPWR _14618_/A sky130_fd_sc_hd__buf_1
X_13706_ _13704_/Y _13705_/Y _13651_/Y VGND VGND VPWR VPWR _13777_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16425_ _16416_/Y _16437_/B _16415_/A VGND VGND VPWR VPWR _16434_/A sky130_fd_sc_hd__a21oi_1
X_14686_ _15349_/A _14742_/B VGND VGND VPWR VPWR _14686_/Y sky130_fd_sc_hd__nand2_1
X_11898_ _12997_/A _11898_/B VGND VGND VPWR VPWR _11898_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13637_ _15125_/A _13637_/B VGND VGND VPWR VPWR _13637_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10849_ _09424_/A _09424_/B _09424_/Y VGND VGND VPWR VPWR _10850_/A sky130_fd_sc_hd__o21ai_1
X_16356_ _08230_/X _16466_/Q _08233_/X _16402_/B _16343_/X VGND VGND VPWR VPWR _16466_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_118_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13568_ _13568_/A VGND VGND VPWR VPWR _13568_/Y sky130_fd_sc_hd__inv_2
X_16287_ _16334_/A _16334_/B VGND VGND VPWR VPWR _16287_/Y sky130_fd_sc_hd__nor2_1
X_12519_ _12519_/A _12519_/B VGND VGND VPWR VPWR _12519_/Y sky130_fd_sc_hd__nand2_1
X_15307_ _15278_/X _15306_/Y _15278_/X _15306_/Y VGND VGND VPWR VPWR _15343_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15238_ _15184_/A _15184_/B _15184_/Y VGND VGND VPWR VPWR _15238_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13499_ _11334_/X _13490_/X _11334_/X _13490_/X VGND VGND VPWR VPWR _13500_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_99_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15169_ _15107_/A _15107_/B _15107_/Y _15099_/X VGND VGND VPWR VPWR _15169_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09730_ _09730_/A _09730_/B VGND VGND VPWR VPWR _09733_/A sky130_fd_sc_hd__or2_1
XFILLER_95_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09661_ _09591_/Y _09659_/X _09660_/Y VGND VGND VPWR VPWR _09661_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08612_ _08612_/A VGND VGND VPWR VPWR _08612_/Y sky130_fd_sc_hd__clkinvlp_2
X_09592_ _09490_/A _09490_/B _09490_/Y VGND VGND VPWR VPWR _09592_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08543_ _08543_/A _08543_/B VGND VGND VPWR VPWR _09860_/A sky130_fd_sc_hd__or2_2
X_08474_ input16/X input32/X VGND VGND VPWR VPWR _08474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09026_ _08645_/X _09007_/Y _08645_/X _09007_/Y VGND VGND VPWR VPWR _09539_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09928_ _09928_/A _09928_/B VGND VGND VPWR VPWR _09928_/X sky130_fd_sc_hd__and2_1
XFILLER_58_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09859_ _09859_/A _09859_/B VGND VGND VPWR VPWR _09914_/A sky130_fd_sc_hd__or2_1
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12870_ _12859_/A _12859_/B _12859_/Y VGND VGND VPWR VPWR _12870_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11821_ _13628_/A _11846_/B VGND VGND VPWR VPWR _11821_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14540_/A _14521_/X VGND VGND VPWR VPWR _14540_/X sky130_fd_sc_hd__or2b_1
XFILLER_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11752_ _11753_/A _11753_/B VGND VGND VPWR VPWR _11752_/X sky130_fd_sc_hd__and2_1
XFILLER_26_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11681_/Y _11682_/X _11681_/Y _11682_/X VGND VGND VPWR VPWR _11683_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10703_ _13636_/A _10791_/B _10702_/Y VGND VGND VPWR VPWR _10703_/Y sky130_fd_sc_hd__o21ai_1
X_14471_ _15038_/A _11917_/Y _11865_/Y _14436_/X VGND VGND VPWR VPWR _14471_/X sky130_fd_sc_hd__o22a_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16210_ _16255_/B VGND VGND VPWR VPWR _16322_/A sky130_fd_sc_hd__clkbuf_2
X_13422_ _14100_/A _13425_/B VGND VGND VPWR VPWR _13422_/Y sky130_fd_sc_hd__nor2_1
X_10634_ _11885_/A VGND VGND VPWR VPWR _12997_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16141_ _16140_/A _16139_/Y _16140_/Y _16139_/A _16388_/A VGND VGND VPWR VPWR _16273_/A
+ sky130_fd_sc_hd__a221o_1
X_13353_ _15473_/A _13354_/B VGND VGND VPWR VPWR _13402_/A sky130_fd_sc_hd__and2_1
XFILLER_10_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12304_ _12248_/X _12303_/Y _12248_/X _12303_/Y VGND VGND VPWR VPWR _12305_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10565_ _10564_/A _10563_/Y _10564_/Y _10563_/A _10976_/A VGND VGND VPWR VPWR _10677_/B
+ sky130_fd_sc_hd__a221o_1
X_16072_ _16041_/X _16071_/Y _16041_/X _16071_/Y VGND VGND VPWR VPWR _16110_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13284_ _13284_/A VGND VGND VPWR VPWR _13284_/Y sky130_fd_sc_hd__inv_2
X_10496_ _13620_/A _10529_/B VGND VGND VPWR VPWR _10496_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12235_ _12235_/A _12136_/X VGND VGND VPWR VPWR _12235_/X sky130_fd_sc_hd__or2b_1
X_15023_ _11740_/Y _14998_/X _11740_/Y _14998_/X VGND VGND VPWR VPWR _15030_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12166_ _12165_/Y _12074_/X _12097_/Y VGND VGND VPWR VPWR _12166_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11117_ _11115_/Y _11116_/Y _10997_/Y VGND VGND VPWR VPWR _11291_/A sky130_fd_sc_hd__o21ai_1
XFILLER_122_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12097_ _12097_/A _12165_/B VGND VGND VPWR VPWR _12097_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15925_ _15898_/A _15898_/B _15898_/Y VGND VGND VPWR VPWR _15925_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11048_ _13567_/A VGND VGND VPWR VPWR _12841_/A sky130_fd_sc_hd__buf_1
Xinput8 wbs_adr_i[15] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__buf_1
X_15856_ _15908_/A _15908_/B VGND VGND VPWR VPWR _15856_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14807_ _14807_/A _14807_/B VGND VGND VPWR VPWR _14807_/X sky130_fd_sc_hd__or2_1
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15787_ _16089_/A _15790_/B VGND VGND VPWR VPWR _15787_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12999_ _12927_/X _12998_/Y _12927_/X _12998_/Y VGND VGND VPWR VPWR _13015_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14738_ _14738_/A _14738_/B VGND VGND VPWR VPWR _14738_/X sky130_fd_sc_hd__or2_1
XFILLER_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14669_ _14599_/A _14599_/B _14592_/X _14599_/Y VGND VGND VPWR VPWR _14669_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16408_ _16399_/Y _16407_/Y _16393_/Y VGND VGND VPWR VPWR _16409_/A sky130_fd_sc_hd__o21ai_1
X_16339_ _16281_/Y _16337_/X _16338_/Y VGND VGND VPWR VPWR _16339_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09713_ _09713_/A VGND VGND VPWR VPWR _09714_/B sky130_fd_sc_hd__inv_2
XFILLER_95_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09644_ _09544_/X _09643_/X _09544_/X _09643_/X VGND VGND VPWR VPWR _10735_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ _09484_/A _09484_/B _09484_/Y VGND VGND VPWR VPWR _09575_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08526_ _08694_/A _10120_/B VGND VGND VPWR VPWR _08871_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08457_ _10009_/A VGND VGND VPWR VPWR _09330_/A sky130_fd_sc_hd__inv_2
XFILLER_51_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08388_ _08388_/A VGND VGND VPWR VPWR _08388_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10350_ _10350_/A _10350_/B VGND VGND VPWR VPWR _10521_/A sky130_fd_sc_hd__or2_1
XFILLER_3_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10281_ _10281_/A VGND VGND VPWR VPWR _10350_/A sky130_fd_sc_hd__inv_2
X_09009_ _08962_/X _09025_/S _08631_/Y VGND VGND VPWR VPWR _09024_/S sky130_fd_sc_hd__o21ai_1
X_12020_ _13196_/A _12063_/B VGND VGND VPWR VPWR _12020_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13971_ _13971_/A VGND VGND VPWR VPWR _13972_/B sky130_fd_sc_hd__inv_2
XFILLER_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15710_ _16055_/A _15696_/B _15696_/Y VGND VGND VPWR VPWR _15710_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12922_ _13005_/A _12922_/B VGND VGND VPWR VPWR _12922_/Y sky130_fd_sc_hd__nor2_1
X_15641_ _15641_/A VGND VGND VPWR VPWR _15641_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12853_ _12853_/A _12853_/B VGND VGND VPWR VPWR _12853_/Y sky130_fd_sc_hd__nand2_1
X_15572_ _15595_/A VGND VGND VPWR VPWR _15700_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12784_/A _12784_/B VGND VGND VPWR VPWR _12784_/Y sky130_fd_sc_hd__nand2_1
X_11804_ _11804_/A VGND VGND VPWR VPWR _11850_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_42_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14523_/A VGND VGND VPWR VPWR _15190_/A sky130_fd_sc_hd__buf_1
X_11735_ _11734_/A _11734_/B _11733_/Y _11734_/Y VGND VGND VPWR VPWR _11745_/B sky130_fd_sc_hd__o2bb2a_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _13274_/A _14428_/B _14428_/Y VGND VGND VPWR VPWR _14454_/X sky130_fd_sc_hd__a21o_1
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13405_ _13405_/A _13405_/B VGND VGND VPWR VPWR _14239_/A sky130_fd_sc_hd__or2_2
X_11666_ _11666_/A VGND VGND VPWR VPWR _11666_/Y sky130_fd_sc_hd__clkinvlp_2
X_14385_ _14385_/A _15956_/A VGND VGND VPWR VPWR _15620_/B sky130_fd_sc_hd__or2_1
X_10617_ _10621_/A _10758_/B VGND VGND VPWR VPWR _11892_/A sky130_fd_sc_hd__or2b_1
X_11597_ _09569_/A _09999_/B _10000_/A VGND VGND VPWR VPWR _11598_/A sky130_fd_sc_hd__o21ai_1
XFILLER_128_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16124_ _16061_/X _16122_/X _16133_/B VGND VGND VPWR VPWR _16124_/X sky130_fd_sc_hd__o21a_1
X_13336_ _13281_/A _13335_/Y _13281_/A _13335_/Y VGND VGND VPWR VPWR _13337_/B sky130_fd_sc_hd__a2bb2o_1
X_10548_ _09981_/A _09981_/B _09981_/Y VGND VGND VPWR VPWR _10549_/A sky130_fd_sc_hd__o21ai_1
X_16055_ _16055_/A _16055_/B VGND VGND VPWR VPWR _16059_/B sky130_fd_sc_hd__or2_1
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13267_ _13183_/X _13266_/Y _13183_/X _13266_/Y VGND VGND VPWR VPWR _13274_/B sky130_fd_sc_hd__a2bb2o_1
X_12218_ _12218_/A _12147_/X VGND VGND VPWR VPWR _12218_/X sky130_fd_sc_hd__or2b_1
X_10479_ _11848_/A _10540_/B _11848_/A _10540_/B VGND VGND VPWR VPWR _10479_/X sky130_fd_sc_hd__a2bb2o_1
X_15006_ _12090_/A _15005_/X _12089_/X VGND VGND VPWR VPWR _15006_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13198_ _13198_/A _13198_/B VGND VGND VPWR VPWR _13198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12149_ _13909_/A _12149_/B VGND VGND VPWR VPWR _12149_/X sky130_fd_sc_hd__or2_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15908_ _15908_/A _15908_/B VGND VGND VPWR VPWR _15908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15839_ _15839_/A _15839_/B VGND VGND VPWR VPWR _15840_/A sky130_fd_sc_hd__or2_1
XFILLER_64_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09360_ _09478_/B _09863_/A _09346_/A VGND VGND VPWR VPWR _09360_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08311_ _08311_/A input21/X VGND VGND VPWR VPWR _08312_/B sky130_fd_sc_hd__nor2_1
X_09291_ _08935_/A _08398_/Y _09234_/A _09628_/A VGND VGND VPWR VPWR _09292_/A sky130_fd_sc_hd__a31o_1
XFILLER_60_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08242_ _08242_/A input6/X VGND VGND VPWR VPWR _08307_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09627_ _09627_/A VGND VGND VPWR VPWR _09707_/A sky130_fd_sc_hd__inv_2
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09558_ _08690_/A _09017_/A _09530_/Y _09557_/X VGND VGND VPWR VPWR _09558_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08509_ _08509_/A VGND VGND VPWR VPWR _08656_/A sky130_fd_sc_hd__inv_2
X_11520_ _11516_/Y _12685_/A _11315_/X _11519_/Y VGND VGND VPWR VPWR _11520_/X sky130_fd_sc_hd__o22a_1
XFILLER_11_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09489_ _08789_/A _09469_/X _08789_/A _09469_/X VGND VGND VPWR VPWR _09490_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11451_ _12351_/A _11455_/B VGND VGND VPWR VPWR _11451_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14170_ _14170_/A _12640_/X VGND VGND VPWR VPWR _14170_/X sky130_fd_sc_hd__or2b_1
X_11382_ _11393_/A _11382_/B VGND VGND VPWR VPWR _12314_/A sky130_fd_sc_hd__or2_1
X_10402_ _10402_/A VGND VGND VPWR VPWR _10402_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13121_ _15240_/A _13121_/B VGND VGND VPWR VPWR _13121_/Y sky130_fd_sc_hd__nand2_1
X_10333_ _11787_/A VGND VGND VPWR VPWR _13529_/A sky130_fd_sc_hd__buf_1
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13052_ _15240_/A _13121_/B VGND VGND VPWR VPWR _13052_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10264_ _11577_/A _10237_/B _10237_/X _11602_/A VGND VGND VPWR VPWR _10264_/Y sky130_fd_sc_hd__a22oi_1
X_12003_ _12778_/A _12078_/A _12002_/Y VGND VGND VPWR VPWR _12003_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10195_ _10122_/Y _10193_/Y _10194_/Y VGND VGND VPWR VPWR _10195_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13954_ _13904_/Y _13952_/X _13953_/Y VGND VGND VPWR VPWR _13954_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13885_ _14832_/A _13990_/B VGND VGND VPWR VPWR _13885_/Y sky130_fd_sc_hd__nand2_1
X_12905_ _12928_/A VGND VGND VPWR VPWR _14460_/A sky130_fd_sc_hd__buf_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _15624_/A VGND VGND VPWR VPWR _15624_/Y sky130_fd_sc_hd__inv_2
X_12836_ _12917_/A VGND VGND VPWR VPWR _12836_/X sky130_fd_sc_hd__buf_1
XFILLER_62_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15488_/Y _15553_/Y _15554_/Y VGND VGND VPWR VPWR _15555_/X sky130_fd_sc_hd__o21a_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _12921_/X _14505_/X _12921_/X _14505_/X VGND VGND VPWR VPWR _14507_/B sky130_fd_sc_hd__a2bb2o_1
X_12767_ _12757_/Y _12765_/X _12766_/Y VGND VGND VPWR VPWR _12767_/X sky130_fd_sc_hd__o21a_1
X_15486_ _14930_/A _15437_/B _15437_/X _15485_/X VGND VGND VPWR VPWR _15486_/X sky130_fd_sc_hd__o22a_1
X_11718_ _11718_/A VGND VGND VPWR VPWR _11791_/A sky130_fd_sc_hd__inv_2
X_12698_ _10381_/A _12661_/A _10381_/Y _12661_/Y VGND VGND VPWR VPWR _12699_/B sky130_fd_sc_hd__o22a_1
XFILLER_30_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput11 wbs_adr_i[3] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11649_ _12445_/A _11650_/B VGND VGND VPWR VPWR _11649_/X sky130_fd_sc_hd__and2_1
X_14437_ _11866_/Y _14436_/X _11866_/Y _14436_/X VGND VGND VPWR VPWR _14438_/B sky130_fd_sc_hd__o2bb2a_1
Xinput22 wbs_dat_i[13] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_2
XFILLER_30_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14368_ _14375_/A _14375_/B VGND VGND VPWR VPWR _14369_/A sky130_fd_sc_hd__or2_2
Xinput33 wbs_dat_i[9] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_4
X_16107_ _16079_/X _16105_/X _16187_/B VGND VGND VPWR VPWR _16107_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13319_ _13368_/A _13368_/B VGND VGND VPWR VPWR _13381_/A sky130_fd_sc_hd__and2_1
XFILLER_6_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14299_ _14308_/A _14299_/B VGND VGND VPWR VPWR _15970_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16038_ _16038_/A _16038_/B VGND VGND VPWR VPWR _16038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08860_ _09498_/A _08825_/A _08827_/Y _08859_/X VGND VGND VPWR VPWR _08860_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08791_ _10129_/A VGND VGND VPWR VPWR _08793_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09412_ _09412_/A _09412_/B VGND VGND VPWR VPWR _09412_/X sky130_fd_sc_hd__or2_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09343_ _09339_/X _09342_/X _09339_/X _09342_/X VGND VGND VPWR VPWR _09343_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_61_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09274_ _09274_/A _09274_/B VGND VGND VPWR VPWR _09274_/X sky130_fd_sc_hd__or2_1
XFILLER_21_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08989_ _08989_/A VGND VGND VPWR VPWR _08989_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10951_ _12942_/A VGND VGND VPWR VPWR _12097_/A sky130_fd_sc_hd__inv_2
XFILLER_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13670_ _15137_/A _13621_/B _13621_/Y VGND VGND VPWR VPWR _13670_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12621_ _12594_/X _12619_/X _14225_/B VGND VGND VPWR VPWR _12621_/X sky130_fd_sc_hd__o21a_1
X_10882_ _12055_/A VGND VGND VPWR VPWR _10886_/A sky130_fd_sc_hd__inv_2
XFILLER_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12552_ _14916_/A _12351_/B _12351_/Y VGND VGND VPWR VPWR _12553_/A sky130_fd_sc_hd__o21ai_1
X_15340_ _15378_/A _15338_/X _15339_/X VGND VGND VPWR VPWR _15340_/X sky130_fd_sc_hd__o21a_1
X_15271_ _15270_/A _15270_/B _11066_/B _15270_/X VGND VGND VPWR VPWR _15271_/X sky130_fd_sc_hd__o22a_1
X_12483_ _15556_/A _12454_/B _12454_/Y _12482_/Y VGND VGND VPWR VPWR _12483_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11503_ _09929_/Y _11502_/X _09928_/X _09931_/B _10794_/X VGND VGND VPWR VPWR _12948_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14222_ _14087_/X _14222_/B VGND VGND VPWR VPWR _14222_/X sky130_fd_sc_hd__and2b_1
X_11434_ _14035_/A _11231_/B _11231_/Y VGND VGND VPWR VPWR _11434_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11365_ _12305_/A _11365_/B VGND VGND VPWR VPWR _11365_/Y sky130_fd_sc_hd__nand2_1
X_14153_ _12429_/A _11618_/A _11619_/Y _13492_/X VGND VGND VPWR VPWR _14153_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_125_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14084_ _14812_/A _14042_/B _14042_/Y VGND VGND VPWR VPWR _14084_/X sky130_fd_sc_hd__a21o_1
X_13104_ _13095_/Y _13102_/X _13103_/Y VGND VGND VPWR VPWR _13104_/X sky130_fd_sc_hd__o21a_1
X_11296_ _12364_/A VGND VGND VPWR VPWR _13792_/A sky130_fd_sc_hd__buf_1
X_10316_ _10367_/A _11760_/A VGND VGND VPWR VPWR _10316_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13035_ _14836_/A _13035_/B VGND VGND VPWR VPWR _13035_/X sky130_fd_sc_hd__or2_1
X_10247_ _10247_/A _10247_/B VGND VGND VPWR VPWR _10247_/X sky130_fd_sc_hd__and2_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10178_ _10108_/A _10177_/Y _10106_/Y VGND VGND VPWR VPWR _10180_/B sky130_fd_sc_hd__o21ai_1
XFILLER_120_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14986_ _14983_/Y _14985_/X _14983_/Y _14985_/X VGND VGND VPWR VPWR _14986_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13937_ _15396_/A _13937_/B VGND VGND VPWR VPWR _13937_/X sky130_fd_sc_hd__and2_1
XFILLER_93_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13868_ _11275_/A _13785_/B _13867_/Y _13782_/X VGND VGND VPWR VPWR _13868_/X sky130_fd_sc_hd__o22a_1
X_15607_ _15679_/A _15679_/B VGND VGND VPWR VPWR _15607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13799_ _14744_/A _13859_/B VGND VGND VPWR VPWR _13799_/Y sky130_fd_sc_hd__nor2_1
X_12819_ _12767_/X _12818_/Y _12767_/X _12818_/Y VGND VGND VPWR VPWR _12843_/B sky130_fd_sc_hd__a2bb2o_1
X_15538_ _15479_/Y _15537_/X _15479_/Y _15537_/X VGND VGND VPWR VPWR _15539_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15469_ _15397_/X _15468_/X _15397_/X _15468_/X VGND VGND VPWR VPWR _15470_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09961_ _09960_/A _09972_/B _09960_/Y VGND VGND VPWR VPWR _09962_/A sky130_fd_sc_hd__o21ai_1
X_08912_ _08970_/A _08970_/B VGND VGND VPWR VPWR _08912_/X sky130_fd_sc_hd__and2_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _09886_/A _09886_/B _09887_/B VGND VGND VPWR VPWR _09918_/A sky130_fd_sc_hd__a21bo_1
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _08843_/A VGND VGND VPWR VPWR _08844_/A sky130_fd_sc_hd__buf_1
XFILLER_85_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08774_ _08773_/A _08739_/A _08773_/Y _08739_/Y VGND VGND VPWR VPWR _09332_/B sky130_fd_sc_hd__o22a_1
XFILLER_38_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09326_ _10241_/A VGND VGND VPWR VPWR _09327_/B sky130_fd_sc_hd__buf_1
X_09257_ _08819_/A _08817_/A _10069_/A _09256_/X VGND VGND VPWR VPWR _09257_/X sky130_fd_sc_hd__o22a_1
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09188_ _09561_/B _09156_/X _09561_/B _09156_/X VGND VGND VPWR VPWR _09189_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11150_ _12270_/A _11316_/B VGND VGND VPWR VPWR _11150_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10101_ _10099_/A _08679_/B _10100_/Y VGND VGND VPWR VPWR _10108_/A sky130_fd_sc_hd__a21oi_2
XFILLER_103_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11081_ _11236_/A _11079_/X _11080_/X VGND VGND VPWR VPWR _11081_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10032_ _09338_/X _10008_/X _10030_/Y VGND VGND VPWR VPWR _10032_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14840_ _12386_/Y _14839_/X _12386_/Y _14839_/X VGND VGND VPWR VPWR _14841_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14771_ _14771_/A _14771_/B VGND VGND VPWR VPWR _14771_/X sky130_fd_sc_hd__or2_1
XFILLER_63_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13722_ _13774_/A _13774_/B VGND VGND VPWR VPWR _13722_/X sky130_fd_sc_hd__and2_1
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11983_ _13636_/A _11983_/B VGND VGND VPWR VPWR _11983_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10934_ _09990_/A _09660_/B _09660_/Y VGND VGND VPWR VPWR _10934_/X sky130_fd_sc_hd__o21a_1
X_16441_ _16416_/Y _16429_/B _16440_/X VGND VGND VPWR VPWR _16441_/Y sky130_fd_sc_hd__o21ai_1
X_13653_ _13704_/A _13652_/Y _13704_/A _13652_/Y VGND VGND VPWR VPWR _13702_/B sky130_fd_sc_hd__a2bb2o_1
X_10865_ _10437_/A _10864_/A _10437_/Y _10864_/Y _10929_/A VGND VGND VPWR VPWR _12059_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16372_ _16322_/A _16322_/B _16322_/Y VGND VGND VPWR VPWR _16372_/Y sky130_fd_sc_hd__o21ai_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12604_ _12601_/Y _12603_/A _12601_/A _12603_/Y _12502_/A VGND VGND VPWR VPWR _12618_/B
+ sky130_fd_sc_hd__o221a_1
X_13584_ _13583_/A _13583_/B _13644_/A VGND VGND VPWR VPWR _13584_/Y sky130_fd_sc_hd__o21ai_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ _12535_/A _12535_/B VGND VGND VPWR VPWR _12535_/Y sky130_fd_sc_hd__nand2_1
X_15323_ _15333_/A _15333_/B VGND VGND VPWR VPWR _15387_/A sky130_fd_sc_hd__and2_1
X_10796_ _12940_/A VGND VGND VPWR VPWR _12007_/A sky130_fd_sc_hd__inv_2
XFILLER_8_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12466_ _13988_/A _12468_/B VGND VGND VPWR VPWR _12466_/X sky130_fd_sc_hd__and2_1
X_15254_ _15221_/X _15253_/Y _15221_/X _15253_/Y VGND VGND VPWR VPWR _15255_/B sky130_fd_sc_hd__a2bb2o_1
X_11417_ _14046_/A _13349_/A VGND VGND VPWR VPWR _13405_/B sky130_fd_sc_hd__or2_1
X_14205_ _14104_/Y _14204_/X _14104_/Y _14204_/X VGND VGND VPWR VPWR _14206_/B sky130_fd_sc_hd__a2bb2oi_1
X_12397_ _12396_/A _12460_/B _12396_/Y VGND VGND VPWR VPWR _12397_/X sky130_fd_sc_hd__o21a_1
X_15185_ _15119_/A _15119_/B _15119_/Y VGND VGND VPWR VPWR _15185_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14136_ _14137_/A _14138_/A VGND VGND VPWR VPWR _14136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11348_ _11285_/X _11347_/Y _11285_/X _11347_/Y VGND VGND VPWR VPWR _11482_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14067_ _14067_/A _14067_/B VGND VGND VPWR VPWR _14146_/B sky130_fd_sc_hd__or2_1
X_11279_ _11279_/A _11279_/B VGND VGND VPWR VPWR _11279_/X sky130_fd_sc_hd__and2_1
X_13018_ _13085_/A _13016_/X _13017_/X VGND VGND VPWR VPWR _13018_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14969_ _14929_/X _14968_/X _14929_/X _14968_/X VGND VGND VPWR VPWR _14996_/A sky130_fd_sc_hd__a2bb2oi_1
XFILLER_75_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08490_ _08331_/A _08257_/B _08474_/Y _08561_/A VGND VGND VPWR VPWR _08549_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09111_ _09538_/B _09031_/B _09032_/B VGND VGND VPWR VPWR _09112_/A sky130_fd_sc_hd__a21bo_1
XFILLER_31_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09042_ _08843_/A _09459_/B _08719_/Y _09064_/A VGND VGND VPWR VPWR _09042_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09944_ _11846_/A VGND VGND VPWR VPWR _13628_/A sky130_fd_sc_hd__buf_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09875_ _09871_/X _08757_/Y _09871_/X _08757_/Y VGND VGND VPWR VPWR _09888_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _09251_/B VGND VGND VPWR VPWR _10125_/A sky130_fd_sc_hd__clkbuf_2
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08757_ _08757_/A VGND VGND VPWR VPWR _08757_/Y sky130_fd_sc_hd__inv_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08688_ _08688_/A _10117_/B VGND VGND VPWR VPWR _08886_/B sky130_fd_sc_hd__and2_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10650_ _09773_/A _09773_/B _09773_/Y VGND VGND VPWR VPWR _10651_/A sky130_fd_sc_hd__o21ai_1
XFILLER_70_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09309_ _10252_/A _09309_/B VGND VGND VPWR VPWR _09309_/Y sky130_fd_sc_hd__nand2_1
X_10581_ _11870_/A _10654_/B VGND VGND VPWR VPWR _10581_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12320_ _14081_/A _12320_/B VGND VGND VPWR VPWR _12321_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12251_ _13202_/A _12251_/B VGND VGND VPWR VPWR _12251_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11202_ _14020_/A VGND VGND VPWR VPWR _14055_/A sky130_fd_sc_hd__buf_1
X_12182_ _12182_/A _12181_/X VGND VGND VPWR VPWR _12182_/X sky130_fd_sc_hd__or2b_1
XFILLER_1_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11133_ _11133_/A VGND VGND VPWR VPWR _11133_/Y sky130_fd_sc_hd__inv_2
X_15941_ _15887_/X _15940_/Y _15887_/X _15940_/Y VGND VGND VPWR VPWR _15950_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11064_ _11064_/A VGND VGND VPWR VPWR _11066_/B sky130_fd_sc_hd__buf_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10015_ _10015_/A _10015_/B VGND VGND VPWR VPWR _10073_/B sky130_fd_sc_hd__nor2_1
X_15872_ _15872_/A VGND VGND VPWR VPWR _15892_/A sky130_fd_sc_hd__inv_2
XFILLER_91_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14823_ _14790_/A _14790_/B _14790_/X _14822_/X VGND VGND VPWR VPWR _14823_/X sky130_fd_sc_hd__o22a_1
XFILLER_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11966_ _11966_/A _11966_/B VGND VGND VPWR VPWR _11966_/X sky130_fd_sc_hd__or2_1
X_14754_ _14754_/A _14754_/B VGND VGND VPWR VPWR _14754_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10917_ _14622_/A _10870_/B _10870_/X _10916_/X VGND VGND VPWR VPWR _10917_/X sky130_fd_sc_hd__o22a_1
X_14685_ _14665_/X _14684_/Y _14665_/X _14684_/Y VGND VGND VPWR VPWR _14742_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13705_ _13705_/A _13705_/B VGND VGND VPWR VPWR _13705_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16424_ _16421_/Y _16447_/B _16447_/A _16415_/A _16420_/X VGND VGND VPWR VPWR _16426_/A
+ sky130_fd_sc_hd__o221a_1
X_11897_ _11897_/A VGND VGND VPWR VPWR _11897_/Y sky130_fd_sc_hd__inv_2
X_13636_ _13636_/A VGND VGND VPWR VPWR _15125_/A sky130_fd_sc_hd__buf_1
X_10848_ _10924_/A _10925_/B VGND VGND VPWR VPWR _11013_/A sky130_fd_sc_hd__and2_1
XFILLER_20_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16355_ _16331_/X _16354_/Y _16331_/X _16354_/Y VGND VGND VPWR VPWR _16402_/B sky130_fd_sc_hd__a2bb2o_1
X_10779_ _11942_/A _10708_/B _10708_/Y _10778_/X VGND VGND VPWR VPWR _10779_/X sky130_fd_sc_hd__a2bb2o_1
X_13567_ _13567_/A _13567_/B VGND VGND VPWR VPWR _13568_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16286_ _16267_/X _16285_/Y _16267_/X _16285_/Y VGND VGND VPWR VPWR _16334_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12518_ _13443_/A _12305_/B _12305_/Y VGND VGND VPWR VPWR _12519_/B sky130_fd_sc_hd__o21a_1
X_15306_ _14585_/A _15249_/B _15249_/Y VGND VGND VPWR VPWR _15306_/Y sky130_fd_sc_hd__o21ai_1
X_13498_ _13500_/A VGND VGND VPWR VPWR _15051_/A sky130_fd_sc_hd__buf_1
X_15237_ _15237_/A _15237_/B VGND VGND VPWR VPWR _15237_/Y sky130_fd_sc_hd__nand2_1
X_12449_ _13972_/A _12449_/B VGND VGND VPWR VPWR _12449_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15168_ _15167_/A _15167_/B _15167_/Y VGND VGND VPWR VPWR _15168_/X sky130_fd_sc_hd__a21o_1
X_14119_ _14119_/A VGND VGND VPWR VPWR _14876_/A sky130_fd_sc_hd__inv_2
XFILLER_87_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15099_ _15054_/A _15054_/B _15054_/Y _15098_/X VGND VGND VPWR VPWR _15099_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09660_ _09990_/A _09660_/B VGND VGND VPWR VPWR _09660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08611_ _08611_/A VGND VGND VPWR VPWR _08611_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09591_ _09990_/A _09660_/B VGND VGND VPWR VPWR _09591_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08542_ _09472_/B VGND VGND VPWR VPWR _08690_/A sky130_fd_sc_hd__buf_1
XFILLER_63_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08473_ input17/X input33/X VGND VGND VPWR VPWR _08473_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09025_ _08632_/X _08962_/X _09025_/S VGND VGND VPWR VPWR _09538_/B sky130_fd_sc_hd__mux2_1
XFILLER_132_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09927_ _11300_/B _09927_/B VGND VGND VPWR VPWR _09928_/B sky130_fd_sc_hd__nand2b_1
XFILLER_131_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09858_ _09858_/A _09904_/A VGND VGND VPWR VPWR _09859_/B sky130_fd_sc_hd__or2_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08809_ _08810_/B VGND VGND VPWR VPWR _08809_/Y sky130_fd_sc_hd__inv_2
X_09789_ _09753_/Y _11496_/A _09788_/X VGND VGND VPWR VPWR _09789_/X sky130_fd_sc_hd__o21a_1
XFILLER_73_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11820_ _11800_/X _11819_/X _11800_/X _11819_/X VGND VGND VPWR VPWR _11846_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11751_ _10310_/A _11750_/A _10310_/Y _11762_/B VGND VGND VPWR VPWR _11753_/B sky130_fd_sc_hd__o22a_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10702_ _11936_/A _10791_/B VGND VGND VPWR VPWR _10702_/Y sky130_fd_sc_hd__nand2_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11649_/X _11653_/X _11651_/B VGND VGND VPWR VPWR _11682_/X sky130_fd_sc_hd__o21a_1
X_14470_ _14438_/A _14438_/B _14435_/X _14438_/Y VGND VGND VPWR VPWR _14470_/X sky130_fd_sc_hd__o2bb2a_1
X_13421_ _13417_/Y _13419_/Y _13420_/Y VGND VGND VPWR VPWR _13425_/B sky130_fd_sc_hd__o21ai_1
X_10633_ _10633_/A VGND VGND VPWR VPWR _10633_/Y sky130_fd_sc_hd__inv_2
X_16140_ _16140_/A VGND VGND VPWR VPWR _16140_/Y sky130_fd_sc_hd__clkinvlp_2
X_13352_ _11415_/X _13351_/X _11415_/X _13351_/X VGND VGND VPWR VPWR _13354_/B sky130_fd_sc_hd__a2bb2o_1
X_10564_ _10564_/A VGND VGND VPWR VPWR _10564_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16071_ _16042_/A _16042_/B _16042_/Y VGND VGND VPWR VPWR _16071_/Y sky130_fd_sc_hd__o21ai_1
X_12303_ _14011_/A _12205_/B _12205_/Y VGND VGND VPWR VPWR _12303_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13283_ _13255_/Y _13281_/Y _13282_/Y VGND VGND VPWR VPWR _13284_/A sky130_fd_sc_hd__o21ai_1
X_10495_ _10433_/X _10494_/X _10433_/X _10494_/X VGND VGND VPWR VPWR _10529_/B sky130_fd_sc_hd__a2bb2o_1
X_15022_ _15032_/A _15032_/B VGND VGND VPWR VPWR _15076_/A sky130_fd_sc_hd__and2_1
XFILLER_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12234_ _12234_/A _12234_/B VGND VGND VPWR VPWR _12234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12165_ _13705_/A _12165_/B VGND VGND VPWR VPWR _12165_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11116_ _11116_/A VGND VGND VPWR VPWR _11116_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12096_ _12076_/X _12095_/X _12076_/X _12095_/X VGND VGND VPWR VPWR _12165_/B sky130_fd_sc_hd__a2bb2o_1
X_15924_ _15962_/A _15962_/B VGND VGND VPWR VPWR _15924_/X sky130_fd_sc_hd__and2_1
X_11047_ _13921_/A _11082_/B VGND VGND VPWR VPWR _11229_/A sky130_fd_sc_hd__and2_1
XFILLER_77_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15855_ _14283_/X _15850_/X _14283_/X _15850_/X VGND VGND VPWR VPWR _15908_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_37_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 wbs_adr_i[1] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_4
X_14806_ _14806_/A _14806_/B VGND VGND VPWR VPWR _14806_/X sky130_fd_sc_hd__and2_1
XFILLER_92_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15786_ _16245_/A _16241_/A _15785_/X VGND VGND VPWR VPWR _15790_/B sky130_fd_sc_hd__o21ai_1
X_12998_ _14460_/A _12928_/B _12928_/Y VGND VGND VPWR VPWR _12998_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14737_ _14784_/A _14735_/X _14736_/X VGND VGND VPWR VPWR _14737_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11949_ _13692_/A _11904_/B _11904_/Y VGND VGND VPWR VPWR _11949_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14668_ _14668_/A VGND VGND VPWR VPWR _15184_/A sky130_fd_sc_hd__buf_1
XFILLER_32_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16407_ _16407_/A _16407_/B _16407_/C _16407_/D VGND VGND VPWR VPWR _16407_/Y sky130_fd_sc_hd__nor4_1
X_13619_ _15140_/A _13605_/B _13605_/Y _13618_/X VGND VGND VPWR VPWR _13619_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16338_ _16338_/A _16338_/B VGND VGND VPWR VPWR _16338_/Y sky130_fd_sc_hd__nand2_1
X_14599_ _14599_/A _14599_/B VGND VGND VPWR VPWR _14599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16269_ _16162_/Y _16267_/X _16268_/Y VGND VGND VPWR VPWR _16269_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09712_ _09686_/A _09686_/B _09689_/A VGND VGND VPWR VPWR _10216_/A sky130_fd_sc_hd__a21bo_1
XFILLER_67_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09643_ _09538_/A _09538_/B _09538_/X VGND VGND VPWR VPWR _09643_/X sky130_fd_sc_hd__o21ba_1
XFILLER_28_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09574_ _09997_/A _09666_/B VGND VGND VPWR VPWR _09574_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08525_ _08524_/A _08459_/Y _08524_/Y _08459_/A VGND VGND VPWR VPWR _10120_/B sky130_fd_sc_hd__o22a_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08456_ _08532_/A VGND VGND VPWR VPWR _10009_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08387_ _08387_/A _08387_/B VGND VGND VPWR VPWR _08388_/A sky130_fd_sc_hd__or2_1
XFILLER_109_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10280_ _11723_/A VGND VGND VPWR VPWR _13478_/A sky130_fd_sc_hd__buf_1
XFILLER_3_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09008_ _09500_/A _09228_/B _09007_/Y VGND VGND VPWR VPWR _09025_/S sky130_fd_sc_hd__o21ai_1
XFILLER_105_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13970_ _13968_/X _13969_/Y _13968_/X _13969_/Y VGND VGND VPWR VPWR _13971_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12921_ _12921_/A VGND VGND VPWR VPWR _12921_/X sky130_fd_sc_hd__buf_1
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15640_ _15640_/A VGND VGND VPWR VPWR _15640_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12852_ _12808_/Y _12850_/X _12851_/Y VGND VGND VPWR VPWR _12852_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15571_ _15571_/A VGND VGND VPWR VPWR _15595_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11803_ _11801_/A _11801_/B _11801_/X _11802_/Y VGND VGND VPWR VPWR _11850_/B sky130_fd_sc_hd__a22o_1
X_12783_ _12733_/Y _12781_/X _12782_/Y VGND VGND VPWR VPWR _12783_/X sky130_fd_sc_hd__o21a_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14540_/A _14520_/X _14521_/X VGND VGND VPWR VPWR _14522_/X sky130_fd_sc_hd__o21a_1
X_11734_ _11734_/A _11734_/B VGND VGND VPWR VPWR _11734_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14453_ _14460_/A _14460_/B VGND VGND VPWR VPWR _14453_/Y sky130_fd_sc_hd__nor2_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11665_ _09196_/Y _09193_/A _09198_/X _09193_/Y VGND VGND VPWR VPWR _11666_/A sky130_fd_sc_hd__o22a_1
X_13404_ _13404_/A _13404_/B VGND VGND VPWR VPWR _13404_/X sky130_fd_sc_hd__and2_1
X_10616_ _08928_/A _10277_/Y _08929_/B _10277_/A VGND VGND VPWR VPWR _10758_/B sky130_fd_sc_hd__o22a_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14384_ _14341_/X _14382_/X _15628_/B VGND VGND VPWR VPWR _14384_/X sky130_fd_sc_hd__o21a_1
X_11596_ _12446_/A VGND VGND VPWR VPWR _12864_/A sky130_fd_sc_hd__inv_2
X_16123_ _16123_/A _16123_/B VGND VGND VPWR VPWR _16133_/B sky130_fd_sc_hd__or2_1
X_13335_ _14728_/A _13282_/B _13282_/Y VGND VGND VPWR VPWR _13335_/Y sky130_fd_sc_hd__o21ai_1
X_10547_ _13518_/A _10546_/B _10546_/X _10442_/X VGND VGND VPWR VPWR _10547_/X sky130_fd_sc_hd__o22a_1
X_16054_ _16062_/A _16052_/Y _16053_/X VGND VGND VPWR VPWR _16054_/X sky130_fd_sc_hd__o21a_1
X_13266_ _15331_/A _13184_/B _13184_/Y VGND VGND VPWR VPWR _13266_/Y sky130_fd_sc_hd__o21ai_1
X_10478_ _10442_/X _10477_/X _10442_/X _10477_/X VGND VGND VPWR VPWR _10540_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12217_ _12217_/A _12217_/B VGND VGND VPWR VPWR _12217_/Y sky130_fd_sc_hd__nand2_1
X_15005_ _11998_/X _15004_/X _12000_/B VGND VGND VPWR VPWR _15005_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13197_ _13159_/Y _13195_/X _13196_/Y VGND VGND VPWR VPWR _13197_/X sky130_fd_sc_hd__o21a_1
X_12148_ _12218_/A _12146_/X _12147_/X VGND VGND VPWR VPWR _12148_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12079_ _12077_/A _12077_/B _12077_/X _12078_/Y VGND VGND VPWR VPWR _12169_/B sky130_fd_sc_hd__a22o_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15907_ _15904_/Y _15905_/X _15906_/Y VGND VGND VPWR VPWR _15907_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15838_ _15838_/A VGND VGND VPWR VPWR _15839_/B sky130_fd_sc_hd__inv_2
XFILLER_52_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15769_ _14905_/X _15768_/X _14905_/X _15768_/X VGND VGND VPWR VPWR _15770_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_64_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09290_ _10230_/A VGND VGND VPWR VPWR _09297_/A sky130_fd_sc_hd__buf_1
X_08310_ _08308_/Y _08309_/A _08308_/A _08309_/Y _08304_/X VGND VGND VPWR VPWR _08521_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08241_ input22/X VGND VGND VPWR VPWR _08242_/A sky130_fd_sc_hd__inv_4
XFILLER_33_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09626_ _08922_/A _09625_/Y _08922_/A _09625_/Y VGND VGND VPWR VPWR _09952_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_28_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09557_ _08688_/A _09019_/A _09532_/Y _09556_/X VGND VGND VPWR VPWR _09557_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09488_ _09488_/A _09488_/B VGND VGND VPWR VPWR _09488_/Y sky130_fd_sc_hd__nor2_1
X_08508_ _08508_/A VGND VGND VPWR VPWR _09345_/B sky130_fd_sc_hd__inv_2
XFILLER_24_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08439_ _08439_/A VGND VGND VPWR VPWR _08439_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11450_ _11445_/Y _12556_/A _11449_/Y VGND VGND VPWR VPWR _11455_/B sky130_fd_sc_hd__o21ai_1
XFILLER_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10401_ _09303_/A _10235_/A _09303_/Y VGND VGND VPWR VPWR _10403_/A sky130_fd_sc_hd__o21ai_1
X_11381_ _08973_/X _11380_/X _08973_/X _11380_/X VGND VGND VPWR VPWR _11382_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13120_ _13057_/Y _13118_/X _13119_/Y VGND VGND VPWR VPWR _13120_/X sky130_fd_sc_hd__o21a_1
X_10332_ _11722_/A VGND VGND VPWR VPWR _11787_/A sky130_fd_sc_hd__buf_1
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13051_ _13030_/X _13050_/X _13030_/X _13050_/X VGND VGND VPWR VPWR _13121_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12002_ _12778_/A _12078_/A VGND VGND VPWR VPWR _12002_/Y sky130_fd_sc_hd__nor2_1
X_10263_ _09370_/B _10238_/B _10238_/X _11536_/A VGND VGND VPWR VPWR _11602_/A sky130_fd_sc_hd__a22o_1
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10194_ _10194_/A _10194_/B VGND VGND VPWR VPWR _10194_/Y sky130_fd_sc_hd__nand2_1
XFILLER_120_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13953_ _15412_/A _13953_/B VGND VGND VPWR VPWR _13953_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13884_ _13861_/X _13883_/X _13861_/X _13883_/X VGND VGND VPWR VPWR _13990_/B sky130_fd_sc_hd__a2bb2o_1
X_12904_ _14462_/A _12930_/B VGND VGND VPWR VPWR _12904_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _14912_/A _15529_/B _15529_/Y VGND VGND VPWR VPWR _15625_/A sky130_fd_sc_hd__o21ai_1
X_12835_ _10422_/A _12831_/X _10426_/A _12834_/Y VGND VGND VPWR VPWR _12837_/B sky130_fd_sc_hd__o22a_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15554_/A _15554_/B VGND VGND VPWR VPWR _15554_/Y sky130_fd_sc_hd__nand2_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _13609_/Y _13615_/A _15146_/A _13615_/Y VGND VGND VPWR VPWR _14505_/X sky130_fd_sc_hd__a22o_1
X_12766_ _12766_/A _12766_/B VGND VGND VPWR VPWR _12766_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15485_ _14774_/A _15440_/B _15440_/X _15484_/X VGND VGND VPWR VPWR _15485_/X sky130_fd_sc_hd__o22a_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11716_/A _11717_/A2 _11716_/Y VGND VGND VPWR VPWR _11719_/A sky130_fd_sc_hd__a21oi_2
X_12697_ _12697_/A _12697_/B VGND VGND VPWR VPWR _12697_/Y sky130_fd_sc_hd__nor2_1
Xinput12 wbs_adr_i[4] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_4
X_11648_ _11645_/X _11647_/Y _11645_/X _11647_/Y VGND VGND VPWR VPWR _11650_/B sky130_fd_sc_hd__a2bb2o_1
X_14436_ _15036_/A _11851_/Y _11816_/Y _14418_/X VGND VGND VPWR VPWR _14436_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14367_ _14367_/A _14367_/B VGND VGND VPWR VPWR _14375_/B sky130_fd_sc_hd__nor2_1
Xinput23 wbs_dat_i[14] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_4
X_11579_ _11579_/A _11579_/B VGND VGND VPWR VPWR _11579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16106_ _16106_/A _16106_/B VGND VGND VPWR VPWR _16187_/B sky130_fd_sc_hd__or2_1
XFILLER_116_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13318_ _13299_/A _13317_/Y _13299_/A _13317_/Y VGND VGND VPWR VPWR _13368_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14298_ _13444_/X _14297_/X _13444_/X _14297_/X VGND VGND VPWR VPWR _14299_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_6_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16037_ _16016_/Y _16035_/X _16036_/Y VGND VGND VPWR VPWR _16037_/X sky130_fd_sc_hd__o21a_1
X_13249_ _13191_/X _13248_/Y _13191_/X _13248_/Y VGND VGND VPWR VPWR _13285_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08790_ _08789_/A _08733_/A _08789_/Y _08733_/Y VGND VGND VPWR VPWR _10129_/A sky130_fd_sc_hd__o22a_1
XFILLER_96_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09411_ _09412_/A _09412_/B VGND VGND VPWR VPWR _10879_/A sky130_fd_sc_hd__and2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09342_ _09146_/X _09341_/B _09146_/X _09341_/X VGND VGND VPWR VPWR _09342_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09273_ _10244_/A VGND VGND VPWR VPWR _09274_/B sky130_fd_sc_hd__buf_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08988_ _08468_/Y _08987_/X _08468_/Y _08987_/X VGND VGND VPWR VPWR _08988_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10950_ _10948_/Y _10949_/Y _10949_/B _09917_/B _10794_/X VGND VGND VPWR VPWR _12942_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10881_ _09285_/Y _10880_/A _09285_/A _10880_/Y _09445_/A VGND VGND VPWR VPWR _12055_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09609_ _09981_/A _09654_/B VGND VGND VPWR VPWR _09609_/Y sky130_fd_sc_hd__nor2_1
X_12620_ _12620_/A _12620_/B VGND VGND VPWR VPWR _14225_/B sky130_fd_sc_hd__or2_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12551_ _12551_/A VGND VGND VPWR VPWR _12551_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15270_ _15270_/A _15270_/B VGND VGND VPWR VPWR _15270_/X sky130_fd_sc_hd__and2_1
X_12482_ _12482_/A VGND VGND VPWR VPWR _12482_/Y sky130_fd_sc_hd__clkinvlp_2
X_11502_ _09928_/A _09928_/B _09928_/X VGND VGND VPWR VPWR _11502_/X sky130_fd_sc_hd__o21ba_1
X_14221_ _15875_/A _14256_/B VGND VGND VPWR VPWR _14221_/Y sky130_fd_sc_hd__nor2_1
X_11433_ _13397_/A _11437_/B VGND VGND VPWR VPWR _11433_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14152_ _14075_/Y _14151_/X _14075_/Y _14151_/X VGND VGND VPWR VPWR _14152_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11364_ _11262_/X _11363_/Y _11262_/X _11363_/Y VGND VGND VPWR VPWR _11365_/B sky130_fd_sc_hd__a2bb2o_1
X_14083_ _14083_/A _14083_/B VGND VGND VPWR VPWR _14083_/X sky130_fd_sc_hd__and2_1
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13103_ _14563_/A _13103_/B VGND VGND VPWR VPWR _13103_/Y sky130_fd_sc_hd__nand2_1
X_10315_ _11760_/A VGND VGND VPWR VPWR _12701_/A sky130_fd_sc_hd__buf_1
XFILLER_3_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11295_ _11593_/A _11295_/B VGND VGND VPWR VPWR _12364_/A sky130_fd_sc_hd__or2_2
XFILLER_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13034_ _13045_/A _13032_/X _13033_/X VGND VGND VPWR VPWR _13034_/X sky130_fd_sc_hd__o21a_1
X_10246_ _10235_/X _10175_/A _10234_/A VGND VGND VPWR VPWR _10247_/B sky130_fd_sc_hd__o21ai_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10177_ _10177_/A _10177_/B VGND VGND VPWR VPWR _10177_/Y sky130_fd_sc_hd__nor2_1
X_14985_ _14929_/X _14984_/Y _14967_/Y VGND VGND VPWR VPWR _14985_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13936_ _13936_/A VGND VGND VPWR VPWR _13936_/X sky130_fd_sc_hd__buf_1
XFILLER_81_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15606_ _14388_/X _15605_/Y _14388_/X _15605_/Y VGND VGND VPWR VPWR _15679_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13867_ _13867_/A VGND VGND VPWR VPWR _13867_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13798_ _13775_/X _13797_/Y _13775_/X _13797_/Y VGND VGND VPWR VPWR _13859_/B sky130_fd_sc_hd__a2bb2o_1
X_12818_ _12768_/A _12768_/B _12768_/Y VGND VGND VPWR VPWR _12818_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15537_ _15455_/A _15455_/B _15455_/A _15455_/B VGND VGND VPWR VPWR _15537_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12699_/A _12699_/B _12699_/Y VGND VGND VPWR VPWR _12749_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15468_ _15468_/A _15398_/X VGND VGND VPWR VPWR _15468_/X sky130_fd_sc_hd__or2b_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14419_ _11817_/Y _14418_/X _11817_/Y _14418_/X VGND VGND VPWR VPWR _14420_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15399_ _15468_/A _15397_/X _15398_/X VGND VGND VPWR VPWR _15399_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09960_ _09960_/A _09972_/B VGND VGND VPWR VPWR _09960_/Y sky130_fd_sc_hd__nand2_1
X_08911_ _08910_/Y _08860_/X _08910_/Y _08860_/X VGND VGND VPWR VPWR _08970_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09887_/A _09887_/B _09888_/B VGND VGND VPWR VPWR _09923_/A sky130_fd_sc_hd__a21bo_1
XFILLER_112_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _10123_/A VGND VGND VPWR VPWR _08842_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08773_/A VGND VGND VPWR VPWR _08773_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09325_ _09324_/X _08888_/Y _09324_/X _08888_/Y VGND VGND VPWR VPWR _10241_/A sky130_fd_sc_hd__o2bb2a_1
X_09256_ _08962_/X _08825_/A _10065_/A _09255_/X VGND VGND VPWR VPWR _09256_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09187_ _09429_/A _09191_/B VGND VGND VPWR VPWR _11667_/A sky130_fd_sc_hd__nor2_1
XFILLER_134_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11080_ _13925_/A _11080_/B VGND VGND VPWR VPWR _11080_/X sky130_fd_sc_hd__or2_1
X_10100_ _10110_/A VGND VGND VPWR VPWR _10100_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10031_ _10008_/A _10008_/B _10008_/X _10030_/Y VGND VGND VPWR VPWR _10031_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14770_ _14771_/A _14771_/B VGND VGND VPWR VPWR _14772_/A sky130_fd_sc_hd__and2_1
XFILLER_17_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13721_ _13703_/X _13720_/Y _13703_/X _13720_/Y VGND VGND VPWR VPWR _13774_/B sky130_fd_sc_hd__a2bb2o_1
X_11982_ _11980_/Y _11981_/Y _11939_/Y VGND VGND VPWR VPWR _12071_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10933_ _10933_/A VGND VGND VPWR VPWR _11590_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16440_ _16412_/Y _16415_/X _16437_/B _16447_/B VGND VGND VPWR VPWR _16440_/X sky130_fd_sc_hd__o22a_1
X_13652_ _15119_/A _13705_/B _13651_/Y VGND VGND VPWR VPWR _13652_/Y sky130_fd_sc_hd__o21ai_1
X_10864_ _10864_/A VGND VGND VPWR VPWR _10864_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16371_ _16357_/X _16462_/Q _16358_/X _16397_/D _16361_/X VGND VGND VPWR VPWR _16462_/D
+ sky130_fd_sc_hd__o221a_2
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12603_ _12603_/A VGND VGND VPWR VPWR _12603_/Y sky130_fd_sc_hd__clkinvlp_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ _13583_/A _13583_/B VGND VGND VPWR VPWR _13644_/A sky130_fd_sc_hd__nand2_1
X_10795_ _09909_/Y _10793_/X _09908_/X _09911_/B _10794_/X VGND VGND VPWR VPWR _12940_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _13439_/A _12311_/B _12311_/Y VGND VGND VPWR VPWR _12535_/B sky130_fd_sc_hd__o21a_1
X_15322_ _15273_/Y _15321_/X _15273_/Y _15321_/X VGND VGND VPWR VPWR _15333_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_12_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15253_ _15199_/A _15199_/B _15199_/Y VGND VGND VPWR VPWR _15253_/Y sky130_fd_sc_hd__o21ai_1
X_12465_ _12461_/X _12464_/Y _12461_/X _12464_/Y VGND VGND VPWR VPWR _12468_/B sky130_fd_sc_hd__a2bb2o_1
X_14204_ _14105_/A _14105_/B _14105_/Y VGND VGND VPWR VPWR _14204_/X sky130_fd_sc_hd__o21a_1
X_11416_ _11413_/A _11413_/B _11247_/X _11415_/X VGND VGND VPWR VPWR _13349_/A sky130_fd_sc_hd__o211a_1
X_12396_ _12396_/A _12460_/B VGND VGND VPWR VPWR _12396_/Y sky130_fd_sc_hd__nand2_1
X_15184_ _15184_/A _15184_/B VGND VGND VPWR VPWR _15184_/Y sky130_fd_sc_hd__nand2_1
X_14135_ _14062_/X _14134_/Y _14062_/X _14134_/Y VGND VGND VPWR VPWR _14138_/A sky130_fd_sc_hd__a2bb2o_1
X_11347_ _12289_/A _11346_/B _11346_/Y VGND VGND VPWR VPWR _11347_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14066_ _14140_/A _14064_/X _14065_/X VGND VGND VPWR VPWR _14066_/X sky130_fd_sc_hd__o21a_1
X_11278_ _11279_/A VGND VGND VPWR VPWR _14663_/A sky130_fd_sc_hd__buf_1
X_13017_ _14492_/A _13017_/B VGND VGND VPWR VPWR _13017_/X sky130_fd_sc_hd__or2_1
XFILLER_67_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10229_ _09541_/B _09292_/B _08402_/X _10228_/Y VGND VGND VPWR VPWR _10230_/B sky130_fd_sc_hd__o22ai_2
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14968_ _14984_/A _14984_/B _14967_/Y VGND VGND VPWR VPWR _14968_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14899_ _14812_/A _14812_/B _14812_/Y VGND VGND VPWR VPWR _14899_/X sky130_fd_sc_hd__a21o_1
X_13919_ _13844_/X _13918_/Y _13844_/X _13918_/Y VGND VGND VPWR VPWR _13945_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09110_ _09717_/A _09113_/B VGND VGND VPWR VPWR _09110_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09041_ _09041_/A _09041_/B VGND VGND VPWR VPWR _09064_/A sky130_fd_sc_hd__or2_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09943_ _12934_/A VGND VGND VPWR VPWR _11846_/A sky130_fd_sc_hd__inv_2
XFILLER_112_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09874_ _08749_/Y _09873_/A _08749_/A _09937_/B VGND VGND VPWR VPWR _09874_/X sky130_fd_sc_hd__a22o_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _08825_/A VGND VGND VPWR VPWR _09251_/B sky130_fd_sc_hd__inv_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08756_ _09448_/A _09478_/B _08708_/Y VGND VGND VPWR VPWR _08757_/A sky130_fd_sc_hd__a21oi_2
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08687_ _09555_/A _08571_/A _08573_/Y _08686_/X VGND VGND VPWR VPWR _08687_/X sky130_fd_sc_hd__o22a_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09308_ _10252_/A _09309_/B VGND VGND VPWR VPWR _09308_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10580_ _10541_/X _10579_/X _10541_/X _10579_/X VGND VGND VPWR VPWR _10654_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09239_ _09458_/B _09690_/A _09227_/X _09238_/X VGND VGND VPWR VPWR _09239_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12250_ _12201_/X _12156_/X _12203_/B VGND VGND VPWR VPWR _12250_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11201_ _13362_/A VGND VGND VPWR VPWR _14020_/A sky130_fd_sc_hd__inv_2
XFILLER_79_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12181_ _12181_/A _12181_/B VGND VGND VPWR VPWR _12181_/X sky130_fd_sc_hd__or2_1
XFILLER_107_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11132_ _09993_/A _09993_/B _09993_/Y VGND VGND VPWR VPWR _11133_/A sky130_fd_sc_hd__o21ai_1
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15940_ _15888_/A _15888_/B _15888_/Y VGND VGND VPWR VPWR _15940_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11063_ _11063_/A _13753_/B VGND VGND VPWR VPWR _11064_/A sky130_fd_sc_hd__or2_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15871_ _15894_/A _15894_/B VGND VGND VPWR VPWR _15871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10014_ _10014_/A _10014_/B VGND VGND VPWR VPWR _10050_/B sky130_fd_sc_hd__nor2_1
X_14822_ _14794_/A _14794_/B _14794_/X _14821_/X VGND VGND VPWR VPWR _14822_/X sky130_fd_sc_hd__o22a_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11965_ _13101_/A _11964_/B _11066_/B _11964_/X VGND VGND VPWR VPWR _11965_/X sky130_fd_sc_hd__o22a_1
X_14753_ _12279_/Y _14752_/X _12279_/Y _14752_/X VGND VGND VPWR VPWR _14754_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10916_ _14626_/A _10878_/B _10878_/X _10915_/X VGND VGND VPWR VPWR _10916_/X sky130_fd_sc_hd__o22a_1
X_14684_ _14745_/A _14745_/B _14683_/Y VGND VGND VPWR VPWR _14684_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13704_ _13704_/A VGND VGND VPWR VPWR _13704_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16423_ _16468_/Q VGND VGND VPWR VPWR _16447_/A sky130_fd_sc_hd__inv_2
X_11896_ _11888_/Y _11894_/X _11895_/Y VGND VGND VPWR VPWR _11897_/A sky130_fd_sc_hd__o21ai_2
XFILLER_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13635_ _13635_/A VGND VGND VPWR VPWR _13635_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10847_ _10779_/X _10846_/Y _10779_/X _10846_/Y VGND VGND VPWR VPWR _10925_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_13_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16354_ _16332_/A _16332_/B _16332_/Y VGND VGND VPWR VPWR _16354_/Y sky130_fd_sc_hd__o21ai_1
X_10778_ _11976_/A _10716_/B _10716_/Y _10777_/X VGND VGND VPWR VPWR _10778_/X sky130_fd_sc_hd__a2bb2o_1
X_13566_ _13531_/X _13565_/Y _13531_/X _13565_/Y VGND VGND VPWR VPWR _13567_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16285_ _16268_/A _16334_/A _16268_/Y VGND VGND VPWR VPWR _16285_/Y sky130_fd_sc_hd__o21ai_1
X_12517_ _12516_/A _12516_/B _12516_/Y _11710_/X VGND VGND VPWR VPWR _12636_/A sky130_fd_sc_hd__o211a_1
X_15305_ _15345_/A _15345_/B VGND VGND VPWR VPWR _15369_/A sky130_fd_sc_hd__and2_1
X_13497_ _15104_/A _13497_/B VGND VGND VPWR VPWR _13497_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15236_ _15227_/X _15235_/Y _15227_/X _15235_/Y VGND VGND VPWR VPWR _15237_/B sky130_fd_sc_hd__a2bb2o_1
X_12448_ _12443_/X _12447_/X _12443_/X _12447_/X VGND VGND VPWR VPWR _12449_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15167_ _15167_/A _15167_/B VGND VGND VPWR VPWR _15167_/Y sky130_fd_sc_hd__nor2_1
X_12379_ _11521_/A _12272_/Y _12378_/Y VGND VGND VPWR VPWR _12379_/X sky130_fd_sc_hd__a21o_1
X_14118_ _14119_/A _14120_/A VGND VGND VPWR VPWR _14118_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15098_ _15057_/A _15057_/B _15057_/Y _15097_/X VGND VGND VPWR VPWR _15098_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14049_ _14812_/A _14042_/B _14042_/Y _14048_/X VGND VGND VPWR VPWR _14049_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_101_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08610_ _08610_/A _10113_/B VGND VGND VPWR VPWR _08611_/A sky130_fd_sc_hd__or2_1
XFILLER_95_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09590_ _09556_/X _09589_/X _09556_/X _09589_/X VGND VGND VPWR VPWR _09660_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08541_ _09529_/A VGND VGND VPWR VPWR _09472_/B sky130_fd_sc_hd__inv_2
X_08472_ input3/X input19/X VGND VGND VPWR VPWR _08472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09024_ _08819_/A _08618_/X _09024_/S VGND VGND VPWR VPWR _09547_/B sky130_fd_sc_hd__mux2_1
XFILLER_132_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09926_ _11300_/A _11299_/A VGND VGND VPWR VPWR _09927_/B sky130_fd_sc_hd__or2_1
XFILLER_85_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09857_ _09857_/A _09857_/B VGND VGND VPWR VPWR _09904_/A sky130_fd_sc_hd__or2_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08808_ _10127_/A VGND VGND VPWR VPWR _08810_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09788_ _09788_/A _09788_/B VGND VGND VPWR VPWR _09788_/X sky130_fd_sc_hd__or2_1
XFILLER_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08739_ _08739_/A VGND VGND VPWR VPWR _08739_/Y sky130_fd_sc_hd__inv_2
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11750_ _11750_/A VGND VGND VPWR VPWR _11762_/B sky130_fd_sc_hd__inv_2
XFILLER_14_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10701_ _10662_/X _10700_/X _10662_/X _10700_/X VGND VGND VPWR VPWR _10791_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11655_/X _11583_/X _11658_/B VGND VGND VPWR VPWR _11681_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_81_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13420_ _14095_/A _13420_/B VGND VGND VPWR VPWR _13420_/Y sky130_fd_sc_hd__nand2_1
X_10632_ _10615_/Y _10630_/X _10631_/Y VGND VGND VPWR VPWR _10633_/A sky130_fd_sc_hd__o21ai_2
XFILLER_41_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13351_ _14721_/A _13272_/B _13272_/Y VGND VGND VPWR VPWR _13351_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10563_ _10563_/A VGND VGND VPWR VPWR _10563_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16070_ _16112_/A _16112_/B VGND VGND VPWR VPWR _16070_/X sky130_fd_sc_hd__and2_1
X_12302_ _12302_/A _12302_/B VGND VGND VPWR VPWR _12302_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13282_ _14728_/A _13282_/B VGND VGND VPWR VPWR _13282_/Y sky130_fd_sc_hd__nand2_1
X_10494_ _11778_/A _10400_/B _11778_/A _10400_/B VGND VGND VPWR VPWR _10494_/X sky130_fd_sc_hd__a2bb2o_1
X_15021_ _11754_/Y _14999_/X _11754_/Y _14999_/X VGND VGND VPWR VPWR _15032_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12233_ _14047_/A VGND VGND VPWR VPWR _13350_/A sky130_fd_sc_hd__inv_2
X_12164_ _12162_/Y _12163_/Y _12100_/Y VGND VGND VPWR VPWR _12257_/A sky130_fd_sc_hd__o21ai_1
XFILLER_123_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11115_ _12162_/A _11115_/B VGND VGND VPWR VPWR _11115_/Y sky130_fd_sc_hd__nor2_1
X_12095_ _09395_/A _12167_/B _09395_/A _12167_/B VGND VGND VPWR VPWR _12095_/X sky130_fd_sc_hd__a2bb2o_1
X_15923_ _15899_/X _15922_/Y _15899_/X _15922_/Y VGND VGND VPWR VPWR _15962_/B sky130_fd_sc_hd__a2bb2o_1
X_11046_ _10914_/X _11045_/X _10914_/X _11045_/X VGND VGND VPWR VPWR _11082_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15854_ _12650_/Y _15853_/Y _14162_/B VGND VGND VPWR VPWR _15854_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15785_ _15785_/A _15785_/B VGND VGND VPWR VPWR _15785_/X sky130_fd_sc_hd__or2_1
X_14805_ _14725_/Y _14804_/X _14725_/Y _14804_/X VGND VGND VPWR VPWR _14806_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14736_ _14736_/A _14736_/B VGND VGND VPWR VPWR _14736_/X sky130_fd_sc_hd__or2_1
X_12997_ _12997_/A VGND VGND VPWR VPWR _13014_/A sky130_fd_sc_hd__inv_2
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11948_ _11974_/A _11974_/B VGND VGND VPWR VPWR _11948_/Y sky130_fd_sc_hd__nor2_1
X_14667_ _14590_/X _14604_/A _14603_/X VGND VGND VPWR VPWR _14667_/X sky130_fd_sc_hd__o21a_1
X_11879_ _11904_/A _11904_/B VGND VGND VPWR VPWR _11879_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16406_ _16406_/A VGND VGND VPWR VPWR _16406_/Y sky130_fd_sc_hd__inv_2
X_14598_ _14593_/X _14597_/X _14593_/X _14597_/X VGND VGND VPWR VPWR _14599_/B sky130_fd_sc_hd__a2bb2o_1
X_13618_ _12925_/A _13608_/B _13608_/X _13617_/X VGND VGND VPWR VPWR _13618_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16337_ _16284_/Y _16335_/X _16336_/Y VGND VGND VPWR VPWR _16337_/X sky130_fd_sc_hd__o21a_1
X_13549_ _15038_/A _13515_/B _13515_/Y VGND VGND VPWR VPWR _13549_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16268_ _16268_/A _16268_/B VGND VGND VPWR VPWR _16268_/Y sky130_fd_sc_hd__nand2_1
X_16199_ _16104_/A _16104_/B _16104_/Y VGND VGND VPWR VPWR _16199_/X sky130_fd_sc_hd__o21a_1
X_15219_ _15208_/A _15208_/B _15208_/Y _15218_/X VGND VGND VPWR VPWR _15219_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09711_ _09709_/A _09709_/B _09709_/Y _09954_/A VGND VGND VPWR VPWR _09713_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09642_ _09960_/A _09645_/B VGND VGND VPWR VPWR _09642_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09573_ _09559_/X _09572_/X _09559_/X _09572_/X VGND VGND VPWR VPWR _09666_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08524_/A VGND VGND VPWR VPWR _08524_/Y sky130_fd_sc_hd__inv_4
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08455_ _08455_/A1 _08313_/Y _08454_/Y _08313_/A _08441_/X VGND VGND VPWR VPWR _08532_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08386_ _09228_/B VGND VGND VPWR VPWR _08386_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09007_ _08844_/A _09005_/Y _09006_/Y VGND VGND VPWR VPWR _09007_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_117_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09909_ _09734_/A _09904_/Y _09859_/B VGND VGND VPWR VPWR _09909_/Y sky130_fd_sc_hd__o21ai_1
X_12920_ _12920_/A VGND VGND VPWR VPWR _12921_/A sky130_fd_sc_hd__inv_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12851_ _12851_/A _12851_/B VGND VGND VPWR VPWR _12851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11802_ _11802_/A VGND VGND VPWR VPWR _11802_/Y sky130_fd_sc_hd__inv_2
X_15570_ _15655_/B VGND VGND VPWR VPWR _15571_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12782_ _12782_/A _12782_/B VGND VGND VPWR VPWR _12782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _15193_/A _14521_/B VGND VGND VPWR VPWR _14521_/X sky130_fd_sc_hd__or2_1
X_11733_ _11733_/A VGND VGND VPWR VPWR _11733_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11662_/Y _11688_/A _11662_/Y _11688_/A VGND VGND VPWR VPWR _11671_/A sky130_fd_sc_hd__o2bb2a_1
X_14452_ _14431_/X _14451_/X _14431_/X _14451_/X VGND VGND VPWR VPWR _14460_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13403_ _13349_/Y _13402_/X _13349_/Y _13402_/X VGND VGND VPWR VPWR _13404_/B sky130_fd_sc_hd__a2bb2o_1
X_10615_ _11895_/A _10631_/B VGND VGND VPWR VPWR _10615_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16122_ _16138_/A _16140_/A _16121_/X VGND VGND VPWR VPWR _16122_/X sky130_fd_sc_hd__o21a_1
X_14383_ _14383_/A _15954_/A VGND VGND VPWR VPWR _15628_/B sky130_fd_sc_hd__or2_1
XFILLER_6_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11595_ _11595_/A _11595_/B VGND VGND VPWR VPWR _12446_/A sky130_fd_sc_hd__or2_2
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13334_ _13334_/A _13334_/B VGND VGND VPWR VPWR _13334_/X sky130_fd_sc_hd__and2_1
X_10546_ _11804_/A _10546_/B VGND VGND VPWR VPWR _10546_/X sky130_fd_sc_hd__and2_1
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16053_ _16053_/A _16053_/B VGND VGND VPWR VPWR _16053_/X sky130_fd_sc_hd__or2_1
X_13265_ _14428_/A VGND VGND VPWR VPWR _13274_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10477_ _13518_/A _10546_/B _13518_/A _10546_/B VGND VGND VPWR VPWR _10477_/X sky130_fd_sc_hd__a2bb2o_1
X_12216_ _12148_/X _12215_/X _12148_/X _12215_/X VGND VGND VPWR VPWR _12217_/B sky130_fd_sc_hd__a2bb2o_1
X_15004_ _11927_/X _15003_/X _11929_/B VGND VGND VPWR VPWR _15004_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13196_ _13196_/A _13196_/B VGND VGND VPWR VPWR _13196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12147_ _13913_/A _12147_/B VGND VGND VPWR VPWR _12147_/X sky130_fd_sc_hd__or2_1
XFILLER_2_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12078_ _12078_/A VGND VGND VPWR VPWR _12078_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15906_ _15906_/A _15906_/B VGND VGND VPWR VPWR _15906_/Y sky130_fd_sc_hd__nand2_1
X_11029_ _13909_/A _11088_/B VGND VGND VPWR VPWR _11211_/A sky130_fd_sc_hd__and2_1
XFILLER_64_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15837_ _16136_/A VGND VGND VPWR VPWR _16277_/A sky130_fd_sc_hd__inv_2
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15768_ _14906_/A _14906_/B _14906_/Y VGND VGND VPWR VPWR _15768_/X sky130_fd_sc_hd__o21a_1
X_15699_ _15553_/Y _15698_/X _15553_/Y _15698_/X VGND VGND VPWR VPWR _15700_/B sky130_fd_sc_hd__a2bb2oi_1
X_14719_ _11067_/B _14718_/X _11067_/B _14718_/X VGND VGND VPWR VPWR _14721_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08240_ input6/X VGND VGND VPWR VPWR _08306_/B sky130_fd_sc_hd__inv_2
XFILLER_20_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09625_ _09503_/A _09505_/Y _09503_/Y VGND VGND VPWR VPWR _09625_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09556_ _09595_/A _09554_/X _09595_/B VGND VGND VPWR VPWR _09556_/X sky130_fd_sc_hd__o21ba_1
X_09487_ _08781_/A _09471_/X _08781_/A _09471_/X VGND VGND VPWR VPWR _09488_/B sky130_fd_sc_hd__o2bb2a_1
X_08507_ _08507_/A _09677_/B VGND VGND VPWR VPWR _08509_/A sky130_fd_sc_hd__or2_4
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08438_ _08565_/B _08433_/X _09452_/A VGND VGND VPWR VPWR _08439_/A sky130_fd_sc_hd__o21ai_1
XFILLER_24_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08369_ _08266_/A input13/X _08347_/B _08368_/X VGND VGND VPWR VPWR _08418_/A sky130_fd_sc_hd__o22a_1
XFILLER_11_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10400_ _11778_/A _10400_/B VGND VGND VPWR VPWR _10400_/X sky130_fd_sc_hd__and2_1
X_11380_ _08901_/X _11380_/B VGND VGND VPWR VPWR _11380_/X sky130_fd_sc_hd__and2b_1
X_10331_ _09954_/A _10330_/A _09954_/Y _10330_/Y _10445_/A VGND VGND VPWR VPWR _11722_/A
+ sky130_fd_sc_hd__o221a_1
X_13050_ _13050_/A _13031_/X VGND VGND VPWR VPWR _13050_/X sky130_fd_sc_hd__or2b_1
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10262_ _09376_/B _10239_/B _10239_/X _11331_/A VGND VGND VPWR VPWR _11536_/A sky130_fd_sc_hd__a22o_1
XFILLER_127_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12001_ _12082_/B _12000_/Y _12082_/B _12000_/Y VGND VGND VPWR VPWR _12078_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10193_ _10194_/A _10194_/B VGND VGND VPWR VPWR _10193_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13952_ _13908_/Y _13950_/X _13951_/Y VGND VGND VPWR VPWR _13952_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12903_ _12842_/X _12902_/Y _12842_/X _12902_/Y VGND VGND VPWR VPWR _12930_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13883_ _13883_/A _13882_/X VGND VGND VPWR VPWR _13883_/X sky130_fd_sc_hd__or2b_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15622_ _15675_/A _15675_/B VGND VGND VPWR VPWR _15622_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12834_ _12833_/A _12833_/B _12833_/Y VGND VGND VPWR VPWR _12834_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15491_/X _15551_/X _15573_/B VGND VGND VPWR VPWR _15553_/Y sky130_fd_sc_hd__o21ai_2
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12765_ _12761_/Y _12763_/Y _12764_/Y VGND VGND VPWR VPWR _12765_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14504_/A VGND VGND VPWR VPWR _15216_/A sky130_fd_sc_hd__buf_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11716_/A _11716_/B VGND VGND VPWR VPWR _11716_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15484_ _14778_/A _15443_/B _15443_/X _15483_/X VGND VGND VPWR VPWR _15484_/X sky130_fd_sc_hd__o22a_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _10466_/A _12663_/A _10466_/Y _12663_/Y VGND VGND VPWR VPWR _12697_/B sky130_fd_sc_hd__o22a_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14435_ _14420_/A _14420_/B _14420_/Y _14434_/X VGND VGND VPWR VPWR _14435_/X sky130_fd_sc_hd__o2bb2a_1
X_11647_ _11646_/Y _11495_/X _11549_/Y VGND VGND VPWR VPWR _11647_/Y sky130_fd_sc_hd__o21ai_1
Xinput13 wbs_adr_i[5] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_1
Xinput24 wbs_dat_i[15] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_2
X_14366_ _14239_/A _14365_/A _14243_/B _14365_/Y VGND VGND VPWR VPWR _14367_/B sky130_fd_sc_hd__o22a_1
X_11578_ _09362_/A _11577_/Y _09364_/X VGND VGND VPWR VPWR _11579_/B sky130_fd_sc_hd__o21a_1
X_16105_ _16101_/Y _16103_/X _16104_/Y VGND VGND VPWR VPWR _16105_/X sky130_fd_sc_hd__o21a_1
X_13317_ _14740_/A _13300_/B _13300_/Y VGND VGND VPWR VPWR _13317_/Y sky130_fd_sc_hd__o21ai_1
X_10529_ _11842_/A _10529_/B VGND VGND VPWR VPWR _10529_/Y sky130_fd_sc_hd__nand2_1
X_16036_ _16036_/A _16036_/B VGND VGND VPWR VPWR _16036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14297_ _13445_/A _13445_/B _13445_/Y VGND VGND VPWR VPWR _14297_/X sky130_fd_sc_hd__o21a_1
X_13248_ _13192_/A _13192_/B _13192_/Y VGND VGND VPWR VPWR _13248_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13179_ _13832_/A VGND VGND VPWR VPWR _15329_/A sky130_fd_sc_hd__buf_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09410_ _09409_/A _09409_/B _10402_/A _09409_/Y VGND VGND VPWR VPWR _09412_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09341_ _09341_/A _09341_/B VGND VGND VPWR VPWR _09341_/X sky130_fd_sc_hd__and2_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09272_ _09257_/X _08905_/Y _09257_/X _08905_/Y VGND VGND VPWR VPWR _10244_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08987_ _08870_/Y _08985_/X _08986_/Y VGND VGND VPWR VPWR _08987_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10880_ _10880_/A VGND VGND VPWR VPWR _10880_/Y sky130_fd_sc_hd__inv_2
X_09608_ _09550_/X _09607_/Y _09550_/X _09607_/Y VGND VGND VPWR VPWR _09654_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09539_ _09539_/A _09539_/B VGND VGND VPWR VPWR _09539_/X sky130_fd_sc_hd__or2_1
XFILLER_71_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12550_ _12546_/Y _12549_/Y _12546_/A _12549_/A _11710_/A VGND VGND VPWR VPWR _12628_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12481_ _12478_/Y _12479_/Y _12480_/Y VGND VGND VPWR VPWR _12481_/Y sky130_fd_sc_hd__o21ai_1
X_11501_ _11500_/Y _11298_/X _11340_/Y VGND VGND VPWR VPWR _11501_/X sky130_fd_sc_hd__o21a_1
X_14220_ _12621_/X _14219_/X _12621_/X _14219_/X VGND VGND VPWR VPWR _14256_/B sky130_fd_sc_hd__a2bb2o_1
X_11432_ _12587_/A _12586_/A _11431_/X VGND VGND VPWR VPWR _11437_/B sky130_fd_sc_hd__o21ai_1
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14151_ _14149_/X _14150_/X _14149_/X _14150_/X VGND VGND VPWR VPWR _14151_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11363_ _14061_/A _11179_/B _11179_/Y VGND VGND VPWR VPWR _11363_/Y sky130_fd_sc_hd__o21ai_1
X_13102_ _13096_/X _13100_/Y _13101_/Y VGND VGND VPWR VPWR _13102_/X sky130_fd_sc_hd__o21a_1
X_14082_ _14081_/A _14081_/B _14239_/A _14081_/Y VGND VGND VPWR VPWR _14083_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10314_ _10314_/A1 _10313_/A _10248_/Y _10313_/Y _10471_/A VGND VGND VPWR VPWR _11760_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_3_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11294_ _09995_/B _11293_/X _09995_/B _11293_/X VGND VGND VPWR VPWR _11295_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13033_ _14749_/A _13033_/B VGND VGND VPWR VPWR _13033_/X sky130_fd_sc_hd__or2_1
X_10245_ _10245_/A VGND VGND VPWR VPWR _10247_/A sky130_fd_sc_hd__inv_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10176_ _10123_/A _10123_/B _10124_/B VGND VGND VPWR VPWR _10180_/A sky130_fd_sc_hd__a21bo_1
XFILLER_121_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14984_ _14984_/A _14984_/B VGND VGND VPWR VPWR _14984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13935_ _13935_/A _13935_/B VGND VGND VPWR VPWR _13936_/A sky130_fd_sc_hd__or2_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13866_ _13974_/A VGND VGND VPWR VPWR _15110_/A sky130_fd_sc_hd__buf_1
X_15605_ _14323_/X _15605_/B VGND VGND VPWR VPWR _15605_/Y sky130_fd_sc_hd__nand2b_1
X_12817_ _12845_/A _12845_/B VGND VGND VPWR VPWR _12817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13797_ _13795_/X _13797_/B VGND VGND VPWR VPWR _13797_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15536_ _15540_/A _15540_/B VGND VGND VPWR VPWR _15536_/Y sky130_fd_sc_hd__nor2_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12748_ _12772_/A _12772_/B VGND VGND VPWR VPWR _12748_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15467_ _15467_/A _15467_/B VGND VGND VPWR VPWR _15467_/Y sky130_fd_sc_hd__nand2_1
X_12679_ _11614_/X _12678_/X _11614_/X _12678_/X VGND VGND VPWR VPWR _12680_/B sky130_fd_sc_hd__o2bb2a_1
X_14418_ _15034_/A _11802_/Y _11770_/Y _14417_/X VGND VGND VPWR VPWR _14418_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15398_ _15398_/A _15398_/B VGND VGND VPWR VPWR _15398_/X sky130_fd_sc_hd__or2_1
X_14349_ _14252_/A _14348_/Y _14252_/A _14348_/Y VGND VGND VPWR VPWR _14379_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16019_ _16034_/A _16034_/B VGND VGND VPWR VPWR _16019_/Y sky130_fd_sc_hd__nor2_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _09888_/A _09888_/B _09888_/X VGND VGND VPWR VPWR _09928_/A sky130_fd_sc_hd__a21bo_1
X_08910_ _08819_/A _10126_/A _08819_/Y VGND VGND VPWR VPWR _08910_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08944_/B VGND VGND VPWR VPWR _10123_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08772_ _09331_/A _09474_/B _08710_/Y VGND VGND VPWR VPWR _08773_/A sky130_fd_sc_hd__a21oi_2
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09324_ _08893_/X _08792_/Y _10047_/A _09259_/X VGND VGND VPWR VPWR _09324_/X sky130_fd_sc_hd__o22a_1
X_09255_ _10018_/A _08834_/A _10061_/A _09254_/Y VGND VGND VPWR VPWR _09255_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09186_ _09182_/Y _09184_/Y _09185_/Y VGND VGND VPWR VPWR _09191_/B sky130_fd_sc_hd__o21ai_1
XFILLER_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10030_ _10035_/B _10029_/X _10035_/A VGND VGND VPWR VPWR _10030_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_130_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11981_ _11981_/A VGND VGND VPWR VPWR _11981_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10932_ _12068_/A _10845_/B _10845_/Y _10779_/X VGND VGND VPWR VPWR _10932_/X sky130_fd_sc_hd__a2bb2o_1
X_13720_ _13718_/X _13720_/B VGND VGND VPWR VPWR _13720_/Y sky130_fd_sc_hd__nand2b_1
X_13651_ _15119_/A _13705_/B VGND VGND VPWR VPWR _13651_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10863_ _09418_/A _09418_/B _09418_/Y VGND VGND VPWR VPWR _10864_/A sky130_fd_sc_hd__o21ai_1
X_16370_ _16323_/X _16369_/Y _16323_/X _16369_/Y VGND VGND VPWR VPWR _16397_/D sky130_fd_sc_hd__a2bb2o_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12602_ _15512_/A _12324_/B _12324_/X VGND VGND VPWR VPWR _12603_/A sky130_fd_sc_hd__o21ba_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ _13537_/X _13581_/Y _13537_/X _13581_/Y VGND VGND VPWR VPWR _13583_/B sky130_fd_sc_hd__a2bb2o_1
X_10794_ _10794_/A VGND VGND VPWR VPWR _10794_/X sky130_fd_sc_hd__clkbuf_2
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ _12532_/A _12532_/B _12532_/Y _11710_/A VGND VGND VPWR VPWR _12632_/A sky130_fd_sc_hd__o211a_1
X_15321_ _14575_/A _15264_/B _15264_/Y VGND VGND VPWR VPWR _15321_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15252_ _15252_/A _15252_/B VGND VGND VPWR VPWR _15252_/Y sky130_fd_sc_hd__nand2_1
X_14203_ _15866_/A _14265_/B VGND VGND VPWR VPWR _14203_/Y sky130_fd_sc_hd__nor2_1
X_12464_ _12459_/X _12464_/B VGND VGND VPWR VPWR _12464_/Y sky130_fd_sc_hd__nand2b_1
X_11415_ _13935_/A _12234_/B VGND VGND VPWR VPWR _11415_/X sky130_fd_sc_hd__or2_1
X_12395_ _12366_/X _12394_/Y _12366_/X _12394_/Y VGND VGND VPWR VPWR _12460_/B sky130_fd_sc_hd__a2bb2o_1
X_15183_ _15156_/X _15182_/Y _15156_/X _15182_/Y VGND VGND VPWR VPWR _15184_/B sky130_fd_sc_hd__a2bb2o_1
X_14134_ _14008_/X _14134_/B VGND VGND VPWR VPWR _14134_/Y sky130_fd_sc_hd__nand2b_1
X_11346_ _12289_/A _11346_/B VGND VGND VPWR VPWR _11346_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14065_ _14065_/A _14065_/B VGND VGND VPWR VPWR _14065_/X sky130_fd_sc_hd__or2_1
X_11277_ _15054_/A VGND VGND VPWR VPWR _13889_/A sky130_fd_sc_hd__buf_1
XFILLER_79_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13016_ _13090_/A _13013_/X _13015_/X VGND VGND VPWR VPWR _13016_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10228_ _10228_/A _10228_/B VGND VGND VPWR VPWR _10228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10159_ _10159_/A _10159_/B VGND VGND VPWR VPWR _10159_/Y sky130_fd_sc_hd__nor2_1
X_14967_ _14984_/A _14984_/B VGND VGND VPWR VPWR _14967_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14898_ _14908_/A _14908_/B VGND VGND VPWR VPWR _14898_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13918_ _14626_/A _13845_/B _13845_/Y VGND VGND VPWR VPWR _13918_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13849_ _14618_/A _13849_/B VGND VGND VPWR VPWR _13849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15519_ _15519_/A _15519_/B VGND VGND VPWR VPWR _15519_/X sky130_fd_sc_hd__or2_1
XFILLER_15_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09040_ _09040_/A VGND VGND VPWR VPWR _09040_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09942_ _09806_/Y _09854_/Y _09854_/B _09897_/B _10794_/A VGND VGND VPWR VPWR _12934_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_131_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09873_ _09873_/A VGND VGND VPWR VPWR _09937_/B sky130_fd_sc_hd__inv_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08823_/X _08726_/X _08823_/A _08726_/X VGND VGND VPWR VPWR _08825_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08755_ _08755_/A VGND VGND VPWR VPWR _09478_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08686_ _09553_/A _08584_/A _08586_/Y _08685_/X VGND VGND VPWR VPWR _08686_/X sky130_fd_sc_hd__o22a_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09307_ _09285_/Y _09305_/Y _09306_/Y VGND VGND VPWR VPWR _09309_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09238_ _09539_/A _09687_/A _09230_/Y _09237_/Y VGND VGND VPWR VPWR _09238_/X sky130_fd_sc_hd__o22a_1
XFILLER_126_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09169_ _09169_/A VGND VGND VPWR VPWR _09750_/A sky130_fd_sc_hd__inv_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12180_ _12181_/A _12181_/B VGND VGND VPWR VPWR _12182_/A sky130_fd_sc_hd__and2_1
X_11200_ _09130_/Y _11199_/A _09130_/A _11199_/Y _11220_/B VGND VGND VPWR VPWR _13362_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_134_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11131_ _13506_/A _11130_/B _11130_/X _10956_/X VGND VGND VPWR VPWR _11131_/X sky130_fd_sc_hd__o22a_1
XFILLER_122_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11062_ _11065_/B VGND VGND VPWR VPWR _13753_/B sky130_fd_sc_hd__inv_2
XFILLER_1_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15870_ _14207_/X _15844_/X _14207_/X _15844_/X VGND VGND VPWR VPWR _15894_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10013_ _10013_/A _10013_/B VGND VGND VPWR VPWR _10047_/B sky130_fd_sc_hd__nor2_1
X_14821_ _14798_/A _14798_/B _14798_/X _14820_/X VGND VGND VPWR VPWR _14821_/X sky130_fd_sc_hd__o22a_1
XFILLER_95_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ _13101_/A _11964_/B VGND VGND VPWR VPWR _11964_/X sky130_fd_sc_hd__and2_1
XFILLER_72_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14752_ _15046_/A _12264_/Y _12184_/Y _14671_/X VGND VGND VPWR VPWR _14752_/X sky130_fd_sc_hd__o22a_1
X_10915_ _14630_/A _10886_/B _10886_/X _10914_/X VGND VGND VPWR VPWR _10915_/X sky130_fd_sc_hd__o22a_1
X_14683_ _14745_/A _14745_/B VGND VGND VPWR VPWR _14683_/Y sky130_fd_sc_hd__nand2_1
X_11895_ _11895_/A _11895_/B VGND VGND VPWR VPWR _11895_/Y sky130_fd_sc_hd__nand2_1
X_13703_ _13723_/A _13701_/X _13702_/X VGND VGND VPWR VPWR _13703_/X sky130_fd_sc_hd__o21a_1
XFILLER_17_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16422_ _16474_/Q _16473_/Q VGND VGND VPWR VPWR _16447_/B sky130_fd_sc_hd__or2_2
X_10846_ _12068_/A _10845_/B _10845_/Y VGND VGND VPWR VPWR _10846_/Y sky130_fd_sc_hd__o21ai_1
X_13634_ _13592_/Y _13631_/Y _13633_/Y VGND VGND VPWR VPWR _13635_/A sky130_fd_sc_hd__o21ai_2
XFILLER_32_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16353_ _08230_/X _16467_/Q _08233_/X _16402_/A _16343_/X VGND VGND VPWR VPWR _16467_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15304_ _15279_/X _15303_/Y _15279_/X _15303_/Y VGND VGND VPWR VPWR _15345_/B sky130_fd_sc_hd__a2bb2o_1
X_10777_ _11974_/A _10724_/B _10724_/Y _10776_/X VGND VGND VPWR VPWR _10777_/X sky130_fd_sc_hd__a2bb2o_1
X_13565_ _15030_/A _13527_/B _13527_/Y VGND VGND VPWR VPWR _13565_/Y sky130_fd_sc_hd__o21ai_1
X_16284_ _16336_/A _16336_/B VGND VGND VPWR VPWR _16284_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12516_ _12516_/A _12516_/B VGND VGND VPWR VPWR _12516_/Y sky130_fd_sc_hd__nand2_1
X_13496_ _11539_/X _13491_/X _11539_/X _13491_/X VGND VGND VPWR VPWR _13497_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15235_ _15181_/A _15181_/B _15181_/Y VGND VGND VPWR VPWR _15235_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12447_ _11632_/A _12441_/B _11632_/A _12441_/B VGND VGND VPWR VPWR _12447_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15166_ _15164_/X _15165_/Y _15164_/X _15165_/Y VGND VGND VPWR VPWR _15167_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14117_ _14056_/X _14116_/X _14056_/X _14116_/X VGND VGND VPWR VPWR _14120_/A sky130_fd_sc_hd__a2bb2o_1
X_12378_ _11321_/A _12272_/A _11521_/B VGND VGND VPWR VPWR _12378_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15097_ _15060_/A _15060_/B _15060_/Y _15096_/X VGND VGND VPWR VPWR _15097_/X sky130_fd_sc_hd__a2bb2o_1
X_11329_ _11317_/X _11328_/Y _11317_/X _11328_/Y VGND VGND VPWR VPWR _11519_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14048_ _14815_/A _14047_/B _14046_/X _14047_/Y VGND VGND VPWR VPWR _14048_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15999_ _15921_/X _15999_/B VGND VGND VPWR VPWR _15999_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_94_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08540_ _08701_/A _08540_/B VGND VGND VPWR VPWR _09529_/A sky130_fd_sc_hd__or2_2
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08471_ input4/X input20/X VGND VGND VPWR VPWR _08471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09023_ _08605_/X _08904_/X _09023_/S VGND VGND VPWR VPWR _09549_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09925_ _09861_/A _09861_/B _09924_/Y VGND VGND VPWR VPWR _11299_/A sky130_fd_sc_hd__a21oi_1
XFILLER_105_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09856_ _09856_/A _09856_/B VGND VGND VPWR VPWR _09857_/B sky130_fd_sc_hd__or2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08807_ _08806_/A _08729_/A _08806_/Y _08729_/Y VGND VGND VPWR VPWR _10127_/A sky130_fd_sc_hd__o22a_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09787_ _09788_/A _09788_/B VGND VGND VPWR VPWR _11496_/A sky130_fd_sc_hd__and2_1
XFILLER_100_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08738_ _08711_/Y _08736_/Y _08737_/X VGND VGND VPWR VPWR _08739_/A sky130_fd_sc_hd__o21ai_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08669_ _09541_/B VGND VGND VPWR VPWR _10228_/A sky130_fd_sc_hd__inv_4
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10666_/X _10798_/B _10666_/X _10798_/B VGND VGND VPWR VPWR _10700_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11677_/Y _11679_/X _11677_/Y _11679_/X VGND VGND VPWR VPWR _11680_/X sky130_fd_sc_hd__a2bb2o_2
X_10631_ _11895_/A _10631_/B VGND VGND VPWR VPWR _10631_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13350_ _13350_/A VGND VGND VPWR VPWR _15473_/A sky130_fd_sc_hd__buf_1
XFILLER_10_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10562_ _10244_/B _10163_/B _10163_/Y VGND VGND VPWR VPWR _10563_/A sky130_fd_sc_hd__a21oi_1
XFILLER_127_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12301_ _12249_/X _12300_/Y _12249_/X _12300_/Y VGND VGND VPWR VPWR _12302_/B sky130_fd_sc_hd__a2bb2o_1
X_13281_ _13281_/A VGND VGND VPWR VPWR _13281_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12232_ _12232_/A _12232_/B VGND VGND VPWR VPWR _12232_/Y sky130_fd_sc_hd__nand2_1
X_10493_ _11842_/A VGND VGND VPWR VPWR _13620_/A sky130_fd_sc_hd__buf_1
X_15020_ _15034_/A _15034_/B VGND VGND VPWR VPWR _15073_/A sky130_fd_sc_hd__and2_1
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12163_ _12163_/A VGND VGND VPWR VPWR _12163_/Y sky130_fd_sc_hd__inv_2
X_11114_ _13048_/A VGND VGND VPWR VPWR _12195_/A sky130_fd_sc_hd__buf_1
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12094_ _12169_/B _12093_/Y _12169_/B _12093_/Y VGND VGND VPWR VPWR _12167_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15922_ _15900_/A _15900_/B _15900_/Y VGND VGND VPWR VPWR _15922_/Y sky130_fd_sc_hd__o21ai_1
X_11045_ _10886_/A _10886_/B _10886_/A _10886_/B VGND VGND VPWR VPWR _11045_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15853_ _15853_/A VGND VGND VPWR VPWR _15853_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15784_ _15784_/A _15784_/B VGND VGND VPWR VPWR _16241_/A sky130_fd_sc_hd__or2_1
X_14804_ _14804_/A _14726_/X VGND VGND VPWR VPWR _14804_/X sky130_fd_sc_hd__or2b_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12996_ _14492_/A _13017_/B VGND VGND VPWR VPWR _13085_/A sky130_fd_sc_hd__and2_1
XFILLER_64_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14735_ _14788_/A _14733_/X _14734_/X VGND VGND VPWR VPWR _14735_/X sky130_fd_sc_hd__o21a_1
X_11947_ _11906_/A _11946_/Y _11906_/A _11946_/Y VGND VGND VPWR VPWR _11974_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14666_ _15240_/A VGND VGND VPWR VPWR _14745_/A sky130_fd_sc_hd__buf_1
X_11878_ _11843_/X _11877_/Y _11843_/X _11877_/Y VGND VGND VPWR VPWR _11904_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16405_ _16399_/Y _16400_/Y _16394_/Y _16393_/Y VGND VGND VPWR VPWR _16406_/A sky130_fd_sc_hd__a31o_1
X_13617_ _13609_/Y _13611_/Y _13616_/Y VGND VGND VPWR VPWR _13617_/X sky130_fd_sc_hd__o21a_1
X_14597_ _14596_/A _14596_/B _14596_/Y VGND VGND VPWR VPWR _14597_/X sky130_fd_sc_hd__a21o_1
X_10829_ _10829_/A _10829_/B VGND VGND VPWR VPWR _10829_/Y sky130_fd_sc_hd__nand2_1
X_16336_ _16336_/A _16336_/B VGND VGND VPWR VPWR _16336_/Y sky130_fd_sc_hd__nand2_1
X_13548_ _13548_/A VGND VGND VPWR VPWR _13548_/Y sky130_fd_sc_hd__inv_2
X_16267_ _16170_/Y _16265_/X _16266_/Y VGND VGND VPWR VPWR _16267_/X sky130_fd_sc_hd__o21a_1
X_15218_ _15211_/A _15211_/B _15211_/Y _15217_/X VGND VGND VPWR VPWR _15218_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13479_ _10421_/B _13478_/Y _11716_/A _10286_/B VGND VGND VPWR VPWR _13480_/A sky130_fd_sc_hd__o22a_1
XFILLER_133_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16198_ _16197_/A _16196_/Y _16197_/Y _16196_/A _15832_/A VGND VGND VPWR VPWR _16257_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15149_ _15140_/A _15140_/B _15140_/Y _15148_/X VGND VGND VPWR VPWR _15149_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09710_ _09683_/A _09683_/B _09686_/A VGND VGND VPWR VPWR _09954_/A sky130_fd_sc_hd__a21bo_2
XFILLER_95_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09641_ _09637_/Y _10743_/A _09640_/Y VGND VGND VPWR VPWR _09645_/B sky130_fd_sc_hd__o21ai_1
XFILLER_83_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09572_ _08694_/A _09152_/A _09526_/A VGND VGND VPWR VPWR _09572_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08523_ _09347_/B _09791_/C VGND VGND VPWR VPWR _08524_/A sky130_fd_sc_hd__or2_1
XFILLER_63_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08454_ _08454_/A VGND VGND VPWR VPWR _08454_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08385_ _08365_/Y _08384_/A _08365_/A _08384_/Y _08303_/A VGND VGND VPWR VPWR _09228_/B
+ sky130_fd_sc_hd__o221a_1
X_09006_ _09006_/A VGND VGND VPWR VPWR _09006_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09908_ _09908_/A _09908_/B VGND VGND VPWR VPWR _09908_/X sky130_fd_sc_hd__and2_1
XFILLER_100_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09839_ _09839_/A VGND VGND VPWR VPWR _09839_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12850_ _12811_/Y _12848_/X _12849_/Y VGND VGND VPWR VPWR _12850_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11801_ _11801_/A _11801_/B VGND VGND VPWR VPWR _11801_/X sky130_fd_sc_hd__or2_1
XFILLER_27_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14544_/A _14518_/X _14519_/X VGND VGND VPWR VPWR _14520_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12781_ _12736_/Y _12779_/X _12780_/Y VGND VGND VPWR VPWR _12781_/X sky130_fd_sc_hd__o21a_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A VGND VGND VPWR VPWR _11734_/A sky130_fd_sc_hd__clkinvlp_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11562_/A _11474_/X _11561_/X VGND VGND VPWR VPWR _11688_/A sky130_fd_sc_hd__o21ai_2
X_14451_ _13925_/A _14426_/B _12141_/A _14426_/B VGND VGND VPWR VPWR _14451_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14382_ _14347_/X _14380_/X _15636_/B VGND VGND VPWR VPWR _14382_/X sky130_fd_sc_hd__o21a_1
X_13402_ _13402_/A _13354_/X VGND VGND VPWR VPWR _13402_/X sky130_fd_sc_hd__or2b_1
X_10614_ _10524_/X _10613_/Y _10524_/X _10613_/Y VGND VGND VPWR VPWR _10631_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16121_ _16121_/A _16121_/B VGND VGND VPWR VPWR _16121_/X sky130_fd_sc_hd__or2_1
X_13333_ _13284_/A _13332_/Y _13284_/A _13332_/Y VGND VGND VPWR VPWR _13334_/B sky130_fd_sc_hd__a2bb2o_1
X_11594_ _09864_/X _09933_/X _09864_/X _09933_/X VGND VGND VPWR VPWR _11595_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_10_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10545_ _11023_/A VGND VGND VPWR VPWR _10545_/X sky130_fd_sc_hd__buf_1
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16052_ _16048_/Y _16050_/X _16051_/Y VGND VGND VPWR VPWR _16052_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13264_ _14724_/A _13276_/B VGND VGND VPWR VPWR _13264_/Y sky130_fd_sc_hd__nor2_1
X_10476_ _10451_/X _10475_/X _10451_/X _10475_/X VGND VGND VPWR VPWR _10546_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12215_ _12215_/A _12149_/X VGND VGND VPWR VPWR _12215_/X sky130_fd_sc_hd__or2b_1
X_13195_ _13162_/Y _13193_/X _13194_/Y VGND VGND VPWR VPWR _13195_/X sky130_fd_sc_hd__o21a_1
X_15003_ _11861_/X _15002_/X _11863_/B VGND VGND VPWR VPWR _15003_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12146_ _12221_/A _12144_/X _12145_/X VGND VGND VPWR VPWR _12146_/X sky130_fd_sc_hd__o21a_1
X_12077_ _12077_/A _12077_/B VGND VGND VPWR VPWR _12077_/X sky130_fd_sc_hd__or2_1
X_15905_ _14177_/X _15849_/X _14177_/X _15849_/X VGND VGND VPWR VPWR _15905_/X sky130_fd_sc_hd__a2bb2o_1
X_11028_ _10917_/X _11027_/X _10917_/X _11027_/X VGND VGND VPWR VPWR _11088_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15836_ _16160_/A _15836_/B VGND VGND VPWR VPWR _16136_/A sky130_fd_sc_hd__or2_1
XFILLER_92_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15767_ _16091_/A VGND VGND VPWR VPWR _16094_/A sky130_fd_sc_hd__buf_6
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12979_ _14411_/A _13025_/B VGND VGND VPWR VPWR _13065_/A sky130_fd_sc_hd__and2_1
X_15698_ _14984_/A _15554_/B _15554_/Y VGND VGND VPWR VPWR _15698_/X sky130_fd_sc_hd__o21a_1
X_14718_ _14643_/A _14643_/B _14643_/Y VGND VGND VPWR VPWR _14718_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14649_ _15335_/A _14649_/B VGND VGND VPWR VPWR _14649_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16319_ _16311_/Y _16317_/X _16318_/Y VGND VGND VPWR VPWR _16319_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09624_ _09957_/A VGND VGND VPWR VPWR _09958_/A sky130_fd_sc_hd__buf_1
XFILLER_102_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09555_ _09555_/A _09555_/B VGND VGND VPWR VPWR _09595_/B sky130_fd_sc_hd__and2_1
XFILLER_24_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09486_ _09486_/A _09486_/B VGND VGND VPWR VPWR _09486_/Y sky130_fd_sc_hd__nor2_1
X_08506_ _08508_/A VGND VGND VPWR VPWR _09863_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08437_ _08712_/A VGND VGND VPWR VPWR _09452_/A sky130_fd_sc_hd__buf_1
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08368_ _08269_/A input12/X _08353_/B _08409_/A VGND VGND VPWR VPWR _08368_/X sky130_fd_sc_hd__o22a_1
X_08299_ _08237_/A input23/X _08238_/A _08296_/A VGND VGND VPWR VPWR _08299_/X sky130_fd_sc_hd__o22a_2
XFILLER_125_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10330_ _10330_/A VGND VGND VPWR VPWR _10330_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10261_ _09382_/B _10240_/B _10240_/X _11155_/A VGND VGND VPWR VPWR _11331_/A sky130_fd_sc_hd__a22o_1
XFILLER_105_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12000_ _11998_/X _12000_/B VGND VGND VPWR VPWR _12000_/Y sky130_fd_sc_hd__nand2b_1
X_10192_ _10238_/B _10139_/B _10139_/Y _10191_/X VGND VGND VPWR VPWR _10194_/B sky130_fd_sc_hd__o2bb2ai_2
XFILLER_78_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13951_ _15410_/A _13951_/B VGND VGND VPWR VPWR _13951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12902_ _12843_/A _12843_/B _12843_/Y VGND VGND VPWR VPWR _12902_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13882_ _13882_/A _13882_/B VGND VGND VPWR VPWR _13882_/X sky130_fd_sc_hd__or2_1
XFILLER_47_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _14384_/X _15620_/Y _14384_/X _15620_/Y VGND VGND VPWR VPWR _15675_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12833_ _12833_/A _12833_/B VGND VGND VPWR VPWR _12833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15552_/A _15552_/B VGND VGND VPWR VPWR _15573_/B sky130_fd_sc_hd__or2_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12764_/A _12764_/B VGND VGND VPWR VPWR _12764_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _14782_/A _15446_/B _15446_/X _15482_/X VGND VGND VPWR VPWR _15483_/X sky130_fd_sc_hd__o22a_1
X_14503_ _15211_/A _14509_/B VGND VGND VPWR VPWR _14564_/A sky130_fd_sc_hd__and2_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _10210_/A _10347_/A _10284_/Y _13478_/B _11724_/B VGND VGND VPWR VPWR _11723_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12695_ _12695_/A _12695_/B VGND VGND VPWR VPWR _12695_/Y sky130_fd_sc_hd__nor2_1
X_14434_ _14422_/A _14422_/B _14422_/Y _14433_/X VGND VGND VPWR VPWR _14434_/X sky130_fd_sc_hd__o2bb2a_1
X_11646_ _12955_/A _11646_/B VGND VGND VPWR VPWR _11646_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 wbs_adr_i[6] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14365_ _14365_/A VGND VGND VPWR VPWR _14365_/Y sky130_fd_sc_hd__inv_2
X_11577_ _11577_/A VGND VGND VPWR VPWR _11577_/Y sky130_fd_sc_hd__inv_2
Xinput25 wbs_dat_i[1] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16104_ _16104_/A _16104_/B VGND VGND VPWR VPWR _16104_/Y sky130_fd_sc_hd__nand2_1
X_14296_ _15972_/A _14402_/B VGND VGND VPWR VPWR _14296_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13316_ _13370_/A _13370_/B VGND VGND VPWR VPWR _13378_/A sky130_fd_sc_hd__and2_1
X_10528_ _10505_/Y _10526_/X _10527_/Y VGND VGND VPWR VPWR _10528_/X sky130_fd_sc_hd__o21a_1
X_16035_ _16019_/Y _16033_/X _16034_/Y VGND VGND VPWR VPWR _16035_/X sky130_fd_sc_hd__o21a_1
X_13247_ _14420_/A VGND VGND VPWR VPWR _14730_/A sky130_fd_sc_hd__buf_1
X_10459_ _10468_/A _10167_/B _10167_/Y VGND VGND VPWR VPWR _10460_/A sky130_fd_sc_hd__a21oi_1
XFILLER_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13178_ _15331_/A _13184_/B VGND VGND VPWR VPWR _13178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12129_ _12052_/X _12128_/Y _12052_/X _12128_/Y VGND VGND VPWR VPWR _12141_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15819_ _16121_/A _15819_/B VGND VGND VPWR VPWR _16150_/B sky130_fd_sc_hd__or2_1
XFILLER_65_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09340_ _09340_/A _09340_/B VGND VGND VPWR VPWR _09341_/B sky130_fd_sc_hd__or2_1
XFILLER_61_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09271_ _09271_/A VGND VGND VPWR VPWR _09274_/A sky130_fd_sc_hd__inv_2
XFILLER_60_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08986_ _08986_/A _08986_/B VGND VGND VPWR VPWR _08986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09607_ _09607_/A _09607_/B VGND VGND VPWR VPWR _09607_/Y sky130_fd_sc_hd__nor2_1
X_09538_ _09538_/A _09538_/B VGND VGND VPWR VPWR _09538_/X sky130_fd_sc_hd__and2_1
XFILLER_52_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11500_ _13780_/A _11500_/B VGND VGND VPWR VPWR _11500_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09469_ _10013_/A _08572_/A _09453_/Y _09468_/X VGND VGND VPWR VPWR _09469_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12480_ _13994_/A _12480_/B VGND VGND VPWR VPWR _12480_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11431_ _15519_/A _11431_/B VGND VGND VPWR VPWR _11431_/X sky130_fd_sc_hd__or2_1
X_11362_ _12305_/A VGND VGND VPWR VPWR _14131_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14150_ _13968_/A _13969_/Y _13967_/X VGND VGND VPWR VPWR _14150_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13101_ _13101_/A _13101_/B VGND VGND VPWR VPWR _13101_/Y sky130_fd_sc_hd__nand2_1
X_10313_ _10313_/A VGND VGND VPWR VPWR _10313_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081_ _14081_/A _14081_/B VGND VGND VPWR VPWR _14081_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11293_ _09785_/A _09785_/B _09785_/Y VGND VGND VPWR VPWR _11293_/X sky130_fd_sc_hd__o21a_1
XFILLER_133_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13032_ _13050_/A _13030_/X _13031_/X VGND VGND VPWR VPWR _13032_/X sky130_fd_sc_hd__o21a_1
X_10244_ _10244_/A _10244_/B VGND VGND VPWR VPWR _10244_/X sky130_fd_sc_hd__or2_1
XFILLER_105_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10175_ _10175_/A VGND VGND VPWR VPWR _10175_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14983_ _14931_/X _14982_/Y _14964_/Y VGND VGND VPWR VPWR _14983_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13934_ _10909_/A _13933_/Y _10909_/A _13933_/Y VGND VGND VPWR VPWR _13937_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13865_ _13863_/Y _13864_/Y _13788_/Y VGND VGND VPWR VPWR _13865_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15604_ _16042_/A VGND VGND VPWR VPWR _15679_/A sky130_fd_sc_hd__inv_2
X_12816_ _12769_/X _12815_/Y _12769_/X _12815_/Y VGND VGND VPWR VPWR _12845_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13796_ _13796_/A _13796_/B VGND VGND VPWR VPWR _13797_/B sky130_fd_sc_hd__or2_1
X_15535_ _15531_/Y _15616_/A _15534_/Y VGND VGND VPWR VPWR _15540_/B sky130_fd_sc_hd__o21ai_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12713_/X _12746_/X _12713_/X _12746_/X VGND VGND VPWR VPWR _12772_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15466_ _15399_/X _15465_/X _15399_/X _15465_/X VGND VGND VPWR VPWR _15467_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12678_ _11615_/Y _12677_/Y _11531_/X VGND VGND VPWR VPWR _12678_/X sky130_fd_sc_hd__o21a_1
X_14417_ _15032_/A _11756_/Y _11775_/Y _14416_/X VGND VGND VPWR VPWR _14417_/X sky130_fd_sc_hd__o22a_1
X_11629_ _11629_/A _11629_/B VGND VGND VPWR VPWR _11629_/X sky130_fd_sc_hd__and2_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15397_ _13935_/A _13935_/B _15395_/X _15471_/A VGND VGND VPWR VPWR _15397_/X sky130_fd_sc_hd__a31o_1
XFILLER_11_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14348_ _15878_/A _14253_/B _14253_/Y VGND VGND VPWR VPWR _14348_/Y sky130_fd_sc_hd__o21ai_1
X_14279_ _13445_/A _14138_/A _14136_/Y VGND VGND VPWR VPWR _14279_/Y sky130_fd_sc_hd__a21oi_1
X_16018_ _15951_/X _16017_/Y _15951_/X _16017_/Y VGND VGND VPWR VPWR _16034_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_97_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08839_/Y _08723_/X _08839_/Y _08723_/X VGND VGND VPWR VPWR _08944_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08771_ _09332_/A VGND VGND VPWR VPWR _09486_/A sky130_fd_sc_hd__buf_1
XFILLER_38_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09323_ _09323_/A _10129_/A VGND VGND VPWR VPWR _10047_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09254_ _09459_/A _10123_/A _08944_/X _09300_/A VGND VGND VPWR VPWR _09254_/Y sky130_fd_sc_hd__a22oi_2
X_09185_ _09430_/A _09185_/B VGND VGND VPWR VPWR _09185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08969_ _08965_/Y _11395_/A _08968_/Y VGND VGND VPWR VPWR _08969_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11980_ _11980_/A _11980_/B VGND VGND VPWR VPWR _11980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10931_ _12106_/A VGND VGND VPWR VPWR _11004_/A sky130_fd_sc_hd__inv_2
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10862_ _10918_/A _10919_/B VGND VGND VPWR VPWR _11027_/A sky130_fd_sc_hd__and2_1
X_13650_ _13645_/X _13649_/Y _13645_/X _13649_/Y VGND VGND VPWR VPWR _13705_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A VGND VGND VPWR VPWR _12601_/Y sky130_fd_sc_hd__inv_2
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13581_ _15042_/A _13509_/B _13509_/Y VGND VGND VPWR VPWR _13581_/Y sky130_fd_sc_hd__o21ai_1
X_10793_ _09908_/A _09908_/B _09908_/X VGND VGND VPWR VPWR _10793_/X sky130_fd_sc_hd__o21ba_1
XFILLER_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ _12532_/A _12532_/B VGND VGND VPWR VPWR _12532_/Y sky130_fd_sc_hd__nand2_1
X_15320_ _15335_/A _15335_/B VGND VGND VPWR VPWR _15384_/A sky130_fd_sc_hd__and2_1
XFILLER_8_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15251_ _15222_/X _15250_/Y _15222_/X _15250_/Y VGND VGND VPWR VPWR _15252_/B sky130_fd_sc_hd__a2bb2o_1
X_12463_ _12459_/X _12461_/X _12464_/B VGND VGND VPWR VPWR _12463_/Y sky130_fd_sc_hd__o21ai_1
X_14202_ _12627_/X _14201_/X _12627_/X _14201_/X VGND VGND VPWR VPWR _14265_/B sky130_fd_sc_hd__a2bb2o_1
X_11414_ _12237_/A VGND VGND VPWR VPWR _14046_/A sky130_fd_sc_hd__inv_2
X_12394_ _12393_/A _12456_/B _12393_/Y VGND VGND VPWR VPWR _12394_/Y sky130_fd_sc_hd__o21ai_1
X_15182_ _15116_/A _15116_/B _15116_/Y VGND VGND VPWR VPWR _15182_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14133_ _14127_/X _14130_/Y _14868_/A _14132_/Y VGND VGND VPWR VPWR _14133_/X sky130_fd_sc_hd__o22a_1
X_11345_ _11494_/A _11344_/Y _11494_/A _11344_/Y VGND VGND VPWR VPWR _11346_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14064_ _14008_/X _14062_/X _14134_/B VGND VGND VPWR VPWR _14064_/X sky130_fd_sc_hd__o21a_1
X_11276_ _12859_/A VGND VGND VPWR VPWR _15054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13015_ _14496_/A _13015_/B VGND VGND VPWR VPWR _13015_/X sky130_fd_sc_hd__or2_1
X_10227_ _10309_/B _10226_/X _10309_/B _10226_/X VGND VGND VPWR VPWR _10296_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10158_ _10128_/A _10128_/B _10129_/B VGND VGND VPWR VPWR _10159_/B sky130_fd_sc_hd__a21bo_1
X_14966_ _14931_/X _14965_/Y _14931_/X _14965_/Y VGND VGND VPWR VPWR _14984_/B sky130_fd_sc_hd__a2bb2o_1
X_10089_ _09749_/X _10034_/B _10034_/Y _10088_/X VGND VGND VPWR VPWR _10089_/X sky130_fd_sc_hd__a2bb2o_1
X_13917_ _13917_/A VGND VGND VPWR VPWR _15404_/A sky130_fd_sc_hd__buf_1
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14897_ _14817_/X _14896_/X _14817_/X _14896_/X VGND VGND VPWR VPWR _14908_/B sky130_fd_sc_hd__a2bb2o_1
X_13848_ _13817_/Y _13846_/X _13847_/Y VGND VGND VPWR VPWR _13848_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13779_ _13777_/Y _13778_/Y _13715_/Y VGND VGND VPWR VPWR _13863_/A sky130_fd_sc_hd__o21ai_1
XFILLER_50_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15518_ _15475_/X _15517_/Y _15475_/X _15517_/Y VGND VGND VPWR VPWR _15640_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15449_ _15449_/A _15449_/B VGND VGND VPWR VPWR _15449_/X sky130_fd_sc_hd__and2_1
XFILLER_129_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09941_ _09941_/A VGND VGND VPWR VPWR _10794_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09872_ _09448_/Y _09871_/X _09478_/X VGND VGND VPWR VPWR _09873_/A sky130_fd_sc_hd__o21ai_2
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08823_/A VGND VGND VPWR VPWR _08823_/X sky130_fd_sc_hd__buf_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _09330_/A VGND VGND VPWR VPWR _09482_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _09551_/A _08596_/A _08598_/Y _08684_/X VGND VGND VPWR VPWR _08685_/X sky130_fd_sc_hd__o22a_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09306_ _10245_/A _09306_/B VGND VGND VPWR VPWR _09306_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09237_ _09237_/A VGND VGND VPWR VPWR _09237_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09168_ _10008_/B _09167_/B _09167_/Y VGND VGND VPWR VPWR _09169_/A sky130_fd_sc_hd__a21oi_2
XFILLER_119_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09099_ _09069_/A _09069_/B _09070_/B VGND VGND VPWR VPWR _09709_/A sky130_fd_sc_hd__o21a_1
XFILLER_134_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11130_ _12080_/A _11130_/B VGND VGND VPWR VPWR _11130_/X sky130_fd_sc_hd__and2_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11061_ _11795_/A VGND VGND VPWR VPWR _13935_/A sky130_fd_sc_hd__buf_1
XFILLER_49_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10012_ _10012_/A _10012_/B VGND VGND VPWR VPWR _10044_/B sky130_fd_sc_hd__nor2_1
X_14820_ _14802_/A _14802_/B _14802_/X _14819_/X VGND VGND VPWR VPWR _14820_/X sky130_fd_sc_hd__o22a_1
XFILLER_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11963_ _11961_/X _11962_/Y _11961_/X _11962_/Y VGND VGND VPWR VPWR _11964_/B sky130_fd_sc_hd__a2bb2o_1
X_14751_ _14673_/A _14673_/B _14670_/X _14673_/Y VGND VGND VPWR VPWR _14751_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10914_ _13824_/A _10894_/B _10894_/Y _10913_/X VGND VGND VPWR VPWR _10914_/X sky130_fd_sc_hd__o2bb2a_1
X_14682_ _14667_/X _14681_/X _14667_/X _14681_/X VGND VGND VPWR VPWR _14745_/B sky130_fd_sc_hd__a2bb2o_1
X_11894_ _11961_/A _11892_/Y _11893_/Y VGND VGND VPWR VPWR _11894_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13702_ _13702_/A _13702_/B VGND VGND VPWR VPWR _13702_/X sky130_fd_sc_hd__or2_1
X_16421_ _16465_/Q VGND VGND VPWR VPWR _16421_/Y sky130_fd_sc_hd__inv_2
X_10845_ _12068_/A _10845_/B VGND VGND VPWR VPWR _10845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13633_ _15128_/A _13633_/B VGND VGND VPWR VPWR _13633_/Y sky130_fd_sc_hd__nand2_1
X_16352_ _16333_/X _16351_/Y _16333_/X _16351_/Y VGND VGND VPWR VPWR _16402_/A sky130_fd_sc_hd__a2bb2o_1
X_15303_ _14587_/A _15246_/B _15246_/Y VGND VGND VPWR VPWR _15303_/Y sky130_fd_sc_hd__o21ai_1
X_10776_ _13078_/A _10733_/B _10733_/Y _10775_/X VGND VGND VPWR VPWR _10776_/X sky130_fd_sc_hd__a2bb2o_1
X_13564_ _13564_/A VGND VGND VPWR VPWR _13564_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16283_ _16269_/X _16282_/Y _16269_/X _16282_/Y VGND VGND VPWR VPWR _16336_/B sky130_fd_sc_hd__o2bb2a_1
X_12515_ _13443_/A _11365_/B _11365_/Y VGND VGND VPWR VPWR _12516_/B sky130_fd_sc_hd__o21a_1
X_13495_ _13495_/A VGND VGND VPWR VPWR _15104_/A sky130_fd_sc_hd__buf_1
XFILLER_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15234_ _15234_/A _15234_/B VGND VGND VPWR VPWR _15234_/Y sky130_fd_sc_hd__nand2_1
X_12446_ _12446_/A VGND VGND VPWR VPWR _13972_/A sky130_fd_sc_hd__buf_1
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15165_ _15100_/X _15103_/X _15105_/B VGND VGND VPWR VPWR _15165_/Y sky130_fd_sc_hd__o21ai_1
X_12377_ _12685_/A _12376_/B _12376_/X _12275_/B VGND VGND VPWR VPWR _12420_/B sky130_fd_sc_hd__a22o_1
XFILLER_126_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14116_ _14116_/A _14057_/X VGND VGND VPWR VPWR _14116_/X sky130_fd_sc_hd__or2b_1
X_11328_ _11328_/A VGND VGND VPWR VPWR _11328_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15096_ _15063_/A _15063_/B _15063_/Y _15095_/X VGND VGND VPWR VPWR _15096_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14047_ _14047_/A _14047_/B VGND VGND VPWR VPWR _14047_/Y sky130_fd_sc_hd__nor2_1
X_11259_ _14108_/A _11213_/B _11213_/Y _11258_/X VGND VGND VPWR VPWR _11259_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15998_ _16053_/A _16053_/B VGND VGND VPWR VPWR _16062_/A sky130_fd_sc_hd__and2_1
XFILLER_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14949_ _14949_/A _14948_/X VGND VGND VPWR VPWR _14949_/X sky130_fd_sc_hd__or2b_1
XFILLER_63_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08470_ input5/X input21/X VGND VGND VPWR VPWR _08470_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09022_ _08795_/X _09011_/Y _08592_/Y _09011_/Y VGND VGND VPWR VPWR _09551_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09924_ _09924_/A VGND VGND VPWR VPWR _09924_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09855_ _09855_/A _09855_/B VGND VGND VPWR VPWR _09897_/B sky130_fd_sc_hd__or2_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08806_ _08806_/A VGND VGND VPWR VPWR _08806_/Y sky130_fd_sc_hd__inv_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09786_ _09995_/B _09784_/Y _09785_/Y VGND VGND VPWR VPWR _09788_/B sky130_fd_sc_hd__o21ai_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08737_ _10011_/A _09529_/A VGND VGND VPWR VPWR _08737_/X sky130_fd_sc_hd__or2_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08668_ _08394_/B _08665_/A _08671_/A _08667_/Y VGND VGND VPWR VPWR _09541_/B sky130_fd_sc_hd__o22a_2
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _13004_/A _10629_/B _10766_/A _10629_/Y VGND VGND VPWR VPWR _10630_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08599_ _08599_/A VGND VGND VPWR VPWR _08599_/Y sky130_fd_sc_hd__clkinvlp_2
X_10561_ _10561_/A VGND VGND VPWR VPWR _11923_/A sky130_fd_sc_hd__inv_2
XFILLER_10_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12300_ _14008_/A _12299_/B _12299_/Y VGND VGND VPWR VPWR _12300_/Y sky130_fd_sc_hd__o21ai_1
X_13280_ _13260_/Y _13278_/Y _13279_/Y VGND VGND VPWR VPWR _13281_/A sky130_fd_sc_hd__o21ai_2
X_10492_ _12930_/A VGND VGND VPWR VPWR _11842_/A sky130_fd_sc_hd__inv_2
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12231_ _12138_/X _12230_/X _12138_/X _12230_/X VGND VGND VPWR VPWR _12232_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12162_ _12162_/A _12162_/B VGND VGND VPWR VPWR _12162_/Y sky130_fd_sc_hd__nor2_1
X_12093_ _12780_/A _12170_/A _12092_/Y VGND VGND VPWR VPWR _12093_/Y sky130_fd_sc_hd__a21oi_1
X_11113_ _11590_/A _11113_/B VGND VGND VPWR VPWR _13048_/A sky130_fd_sc_hd__or2_2
X_15921_ _15964_/A _15964_/B VGND VGND VPWR VPWR _15921_/X sky130_fd_sc_hd__and2_1
XFILLER_103_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11044_ _15078_/A VGND VGND VPWR VPWR _13921_/A sky130_fd_sc_hd__buf_1
XFILLER_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15852_ _14170_/A _15851_/X _12640_/X VGND VGND VPWR VPWR _15853_/A sky130_fd_sc_hd__o21ai_2
XFILLER_64_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15783_ _15777_/A _16028_/A _15656_/A _16028_/B VGND VGND VPWR VPWR _15784_/B sky130_fd_sc_hd__a22o_1
X_14803_ _15464_/A VGND VGND VPWR VPWR _14806_/A sky130_fd_sc_hd__buf_1
X_12995_ _12929_/X _12994_/Y _12929_/X _12994_/Y VGND VGND VPWR VPWR _13017_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14734_ _14734_/A _14734_/B VGND VGND VPWR VPWR _14734_/X sky130_fd_sc_hd__or2_1
X_11946_ _13694_/A _11907_/B _11907_/Y VGND VGND VPWR VPWR _11946_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16404_ _16454_/A _16404_/B VGND VGND VPWR VPWR _16473_/D sky130_fd_sc_hd__or2_1
X_14665_ _14588_/X _14664_/Y _14606_/Y VGND VGND VPWR VPWR _14665_/X sky130_fd_sc_hd__o21a_1
X_11877_ _11844_/A _11844_/B _11844_/Y VGND VGND VPWR VPWR _11877_/Y sky130_fd_sc_hd__o21ai_1
X_13616_ _13005_/A _13615_/Y _12920_/A VGND VGND VPWR VPWR _13616_/Y sky130_fd_sc_hd__o21ai_1
X_14596_ _14596_/A _14596_/B VGND VGND VPWR VPWR _14596_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10828_ _09262_/B _10242_/B _10242_/X VGND VGND VPWR VPWR _10829_/B sky130_fd_sc_hd__a21boi_1
X_16335_ _16287_/Y _16333_/X _16334_/Y VGND VGND VPWR VPWR _16335_/X sky130_fd_sc_hd__o21a_1
X_10759_ _13752_/A VGND VGND VPWR VPWR _10768_/A sky130_fd_sc_hd__inv_2
X_13547_ _13547_/A _13547_/B VGND VGND VPWR VPWR _13548_/A sky130_fd_sc_hd__nand2_1
X_16266_ _16266_/A _16266_/B VGND VGND VPWR VPWR _16266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15217_ _15212_/X _15268_/A _15216_/X VGND VGND VPWR VPWR _15217_/X sky130_fd_sc_hd__o21a_1
X_13478_ _13478_/A _13478_/B VGND VGND VPWR VPWR _13478_/Y sky130_fd_sc_hd__nor2_1
X_16197_ _16197_/A VGND VGND VPWR VPWR _16197_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12429_ _12429_/A _12429_/B VGND VGND VPWR VPWR _12429_/X sky130_fd_sc_hd__or2_1
XFILLER_99_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15148_ _15143_/A _15143_/B _15143_/Y _15147_/X VGND VGND VPWR VPWR _15148_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15079_ _15079_/A _15030_/X VGND VGND VPWR VPWR _15079_/X sky130_fd_sc_hd__or2b_1
XFILLER_68_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09640_ _09958_/A _09640_/B VGND VGND VPWR VPWR _09640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09571_ _09516_/X _09570_/X _09516_/X _09570_/X VGND VGND VPWR VPWR _09997_/A sky130_fd_sc_hd__a2bb2o_1
X_08522_ _09862_/A VGND VGND VPWR VPWR _09347_/B sky130_fd_sc_hd__inv_2
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08453_ _08453_/A VGND VGND VPWR VPWR _08453_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08384_ _08384_/A VGND VGND VPWR VPWR _08384_/Y sky130_fd_sc_hd__inv_2
X_09005_ _08935_/A _09005_/A2 _08664_/X VGND VGND VPWR VPWR _09005_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09907_ _10657_/B _09907_/B VGND VGND VPWR VPWR _09908_/B sky130_fd_sc_hd__nand2b_1
XFILLER_59_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09838_ _09838_/A _09838_/B VGND VGND VPWR VPWR _09839_/A sky130_fd_sc_hd__nand2_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _09769_/A VGND VGND VPWR VPWR _09773_/A sky130_fd_sc_hd__inv_2
XFILLER_132_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11800_ _13559_/A _11773_/B _11773_/X _11799_/X VGND VGND VPWR VPWR _11800_/X sky130_fd_sc_hd__o22a_1
XFILLER_39_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12780_ _12780_/A _12780_/B VGND VGND VPWR VPWR _12780_/Y sky130_fd_sc_hd__nand2_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11731_ _11779_/A _11731_/B VGND VGND VPWR VPWR _11731_/X sky130_fd_sc_hd__or2_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11662_/A _11661_/X VGND VGND VPWR VPWR _11662_/Y sky130_fd_sc_hd__nor2b_1
X_14450_ _14462_/A _14462_/B VGND VGND VPWR VPWR _14450_/Y sky130_fd_sc_hd__nor2_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14381_ _14381_/A _15952_/A VGND VGND VPWR VPWR _15636_/B sky130_fd_sc_hd__or2_1
X_13401_ _13404_/A VGND VGND VPWR VPWR _14904_/A sky130_fd_sc_hd__buf_1
X_10613_ _11838_/A _10525_/B _10525_/Y VGND VGND VPWR VPWR _10613_/Y sky130_fd_sc_hd__o21ai_1
X_11593_ _11593_/A _11593_/B VGND VGND VPWR VPWR _12454_/A sky130_fd_sc_hd__or2_2
X_16120_ _16116_/Y _16147_/A _16119_/Y VGND VGND VPWR VPWR _16140_/A sky130_fd_sc_hd__o21ai_2
X_13332_ _14730_/A _13285_/B _13285_/Y VGND VGND VPWR VPWR _13332_/Y sky130_fd_sc_hd__o21ai_1
X_10544_ _10543_/A _10543_/B _10543_/Y _09392_/A VGND VGND VPWR VPWR _11023_/A sky130_fd_sc_hd__o211a_1
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16051_ _16051_/A _16051_/B VGND VGND VPWR VPWR _16051_/Y sky130_fd_sc_hd__nand2_1
X_13263_ _13185_/X _13262_/Y _13185_/X _13262_/Y VGND VGND VPWR VPWR _13276_/B sky130_fd_sc_hd__a2bb2o_1
X_10475_ _10554_/A _12697_/A _10474_/Y VGND VGND VPWR VPWR _10475_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12214_ _14020_/A _12214_/B VGND VGND VPWR VPWR _12214_/Y sky130_fd_sc_hd__nand2_1
X_13194_ _13194_/A _13194_/B VGND VGND VPWR VPWR _13194_/Y sky130_fd_sc_hd__nand2_1
X_15002_ _11812_/X _15001_/X _11814_/B VGND VGND VPWR VPWR _15002_/X sky130_fd_sc_hd__o21a_1
X_12145_ _13917_/A _12145_/B VGND VGND VPWR VPWR _12145_/X sky130_fd_sc_hd__or2_1
XFILLER_77_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12076_ _13583_/A _12075_/B _12075_/X _11986_/X VGND VGND VPWR VPWR _12076_/X sky130_fd_sc_hd__o22a_1
X_15904_ _15906_/A _15906_/B VGND VGND VPWR VPWR _15904_/Y sky130_fd_sc_hd__nor2_1
X_11027_ _11027_/A _10919_/X VGND VGND VPWR VPWR _11027_/X sky130_fd_sc_hd__or2b_1
X_15835_ _15822_/X _15834_/X _15822_/X _15834_/X VGND VGND VPWR VPWR _15836_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15766_ _15766_/A _15766_/B VGND VGND VPWR VPWR _16091_/A sky130_fd_sc_hd__or2_1
X_12978_ _12937_/X _12977_/Y _12937_/X _12977_/Y VGND VGND VPWR VPWR _13025_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15697_ _15578_/Y _15695_/X _15696_/Y VGND VGND VPWR VPWR _15697_/X sky130_fd_sc_hd__o21a_1
X_14717_ _15398_/A _14717_/B VGND VGND VPWR VPWR _14717_/X sky130_fd_sc_hd__and2_1
XFILLER_72_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11929_ _11927_/X _11929_/B VGND VGND VPWR VPWR _11929_/Y sky130_fd_sc_hd__nand2b_1
X_14648_ _14637_/Y _14646_/Y _14647_/Y VGND VGND VPWR VPWR _14648_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16318_ _16318_/A _16318_/B VGND VGND VPWR VPWR _16318_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14579_ _14579_/A _14579_/B VGND VGND VPWR VPWR _14579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16249_ _16249_/A _16249_/B VGND VGND VPWR VPWR _16249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09623_ _09506_/X _09622_/X _09506_/X _09622_/X VGND VGND VPWR VPWR _09957_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09554_ _09601_/A _09552_/X _09601_/B VGND VGND VPWR VPWR _09554_/X sky130_fd_sc_hd__o21ba_1
XFILLER_102_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09485_ _08773_/A _09473_/X _08773_/A _09473_/X VGND VGND VPWR VPWR _09486_/B sky130_fd_sc_hd__o2bb2a_1
X_08505_ _09146_/A _08505_/B VGND VGND VPWR VPWR _08508_/A sky130_fd_sc_hd__or2_1
XFILLER_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08436_ _10012_/A VGND VGND VPWR VPWR _08712_/A sky130_fd_sc_hd__inv_2
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08367_ _08272_/A input11/X _08364_/B _08366_/A VGND VGND VPWR VPWR _08409_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08298_ _08298_/A VGND VGND VPWR VPWR _08298_/X sky130_fd_sc_hd__buf_1
XFILLER_124_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10260_ _09327_/B _10241_/B _10241_/X _10983_/A VGND VGND VPWR VPWR _11155_/A sky130_fd_sc_hd__a22o_1
XFILLER_133_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10191_ _10239_/B _10143_/B _10143_/Y _10190_/X VGND VGND VPWR VPWR _10191_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13950_ _13912_/Y _13948_/X _13949_/Y VGND VGND VPWR VPWR _13950_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12901_ _12930_/A VGND VGND VPWR VPWR _14462_/A sky130_fd_sc_hd__buf_1
XFILLER_47_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _14335_/X _15620_/B VGND VGND VPWR VPWR _15620_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_100_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13881_ _13882_/A _13882_/B VGND VGND VPWR VPWR _13883_/A sky130_fd_sc_hd__and2_1
XFILLER_74_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12832_ _12832_/A VGND VGND VPWR VPWR _12833_/A sky130_fd_sc_hd__buf_1
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15494_/X _15549_/X _15690_/B VGND VGND VPWR VPWR _15551_/X sky130_fd_sc_hd__o21a_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12830_/A _12833_/B _10422_/A VGND VGND VPWR VPWR _12763_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _14786_/A _15449_/B _15449_/X _15481_/X VGND VGND VPWR VPWR _15482_/X sky130_fd_sc_hd__o22a_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14457_/Y _14501_/X _14457_/Y _14501_/X VGND VGND VPWR VPWR _14509_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_70_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11714_ _11714_/A _11714_/B VGND VGND VPWR VPWR _11724_/B sky130_fd_sc_hd__or2_1
XFILLER_15_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14424_/A _14424_/B _14424_/Y _14432_/X VGND VGND VPWR VPWR _14433_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12694_ _10568_/A _12665_/A _10568_/Y _12665_/Y VGND VGND VPWR VPWR _12695_/B sky130_fd_sc_hd__o22a_1
XFILLER_30_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11645_ _12454_/A _11644_/B _11644_/X VGND VGND VPWR VPWR _11645_/X sky130_fd_sc_hd__a21bo_1
Xinput15 wbs_adr_i[7] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_4
X_14364_ _14904_/A _13404_/B _13404_/X VGND VGND VPWR VPWR _14365_/A sky130_fd_sc_hd__o21ba_1
X_11576_ _15437_/A _11564_/B _11564_/Y _11468_/X VGND VGND VPWR VPWR _11576_/Y sky130_fd_sc_hd__a2bb2oi_1
Xinput26 wbs_dat_i[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_4
X_16103_ _16035_/X _16102_/Y _16035_/X _16102_/Y VGND VGND VPWR VPWR _16103_/X sky130_fd_sc_hd__a2bb2o_1
X_14295_ _14286_/X _14294_/Y _14286_/X _14294_/Y VGND VGND VPWR VPWR _14402_/B sky130_fd_sc_hd__a2bb2o_1
X_13315_ _13302_/A _13314_/Y _13302_/A _13314_/Y VGND VGND VPWR VPWR _13370_/B sky130_fd_sc_hd__a2bb2o_1
X_10527_ _11840_/A _10527_/B VGND VGND VPWR VPWR _10527_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16034_ _16034_/A _16034_/B VGND VGND VPWR VPWR _16034_/Y sky130_fd_sc_hd__nand2_1
X_13246_ _15072_/A VGND VGND VPWR VPWR _14420_/A sky130_fd_sc_hd__inv_2
X_10458_ _10458_/A VGND VGND VPWR VPWR _11857_/A sky130_fd_sc_hd__inv_2
XFILLER_97_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13177_ _13102_/X _13176_/Y _13102_/X _13176_/Y VGND VGND VPWR VPWR _13184_/B sky130_fd_sc_hd__a2bb2o_1
X_10389_ _10368_/X _10388_/X _10368_/X _10388_/X VGND VGND VPWR VPWR _10441_/B sky130_fd_sc_hd__a2bb2o_1
X_12128_ _12039_/A _12053_/B _12053_/Y VGND VGND VPWR VPWR _12128_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12059_ _12059_/A _12059_/B VGND VGND VPWR VPWR _12059_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15818_ _15725_/Y _15816_/X _15817_/Y VGND VGND VPWR VPWR _15818_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15749_ _16108_/A _15809_/B VGND VGND VPWR VPWR _15749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09270_ _09241_/X _09269_/X _09241_/X _09269_/X VGND VGND VPWR VPWR _09271_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08985_ _08875_/X _08983_/X _11462_/B VGND VGND VPWR VPWR _08985_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09606_ _09980_/A VGND VGND VPWR VPWR _09981_/A sky130_fd_sc_hd__buf_1
XFILLER_83_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09537_ _09547_/A _09547_/B VGND VGND VPWR VPWR _09648_/A sky130_fd_sc_hd__nor2_1
X_09468_ _09454_/Y _09466_/X _09467_/X VGND VGND VPWR VPWR _09468_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08419_ _08419_/A VGND VGND VPWR VPWR _08441_/A sky130_fd_sc_hd__clkbuf_2
X_09399_ _09717_/A VGND VGND VPWR VPWR _09412_/A sky130_fd_sc_hd__inv_2
X_11430_ _11254_/X _11429_/Y _11254_/X _11429_/Y VGND VGND VPWR VPWR _12586_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11361_ _11572_/A _11361_/B VGND VGND VPWR VPWR _12305_/A sky130_fd_sc_hd__or2_1
XFILLER_20_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13100_ _14567_/A _13101_/B VGND VGND VPWR VPWR _13100_/Y sky130_fd_sc_hd__nor2_1
X_10312_ _10247_/A _10247_/B _10247_/X VGND VGND VPWR VPWR _10313_/A sky130_fd_sc_hd__o21ba_1
X_14080_ _14046_/X _14079_/X _14046_/A _14079_/X VGND VGND VPWR VPWR _14081_/B sky130_fd_sc_hd__a2bb2o_1
X_11292_ _11290_/Y _11291_/Y _11167_/Y VGND VGND VPWR VPWR _11494_/A sky130_fd_sc_hd__o21ai_1
XFILLER_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13031_ _14668_/A _13031_/B VGND VGND VPWR VPWR _13031_/X sky130_fd_sc_hd__or2_1
X_10243_ _10243_/A _10243_/B VGND VGND VPWR VPWR _10243_/X sky130_fd_sc_hd__or2_1
XFILLER_133_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10174_ _10100_/Y _08647_/A _10111_/A VGND VGND VPWR VPWR _10175_/A sky130_fd_sc_hd__o21ai_2
XFILLER_121_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14982_ _15563_/A _14982_/B VGND VGND VPWR VPWR _14982_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13933_ _14643_/A _13837_/B _13837_/Y VGND VGND VPWR VPWR _13933_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13864_ _15113_/A _13864_/B VGND VGND VPWR VPWR _13864_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15603_ _15602_/A _15601_/Y _15602_/Y _15601_/A _15595_/A VGND VGND VPWR VPWR _16042_/A
+ sky130_fd_sc_hd__a221o_1
X_12815_ _12770_/A _12770_/B _12770_/Y VGND VGND VPWR VPWR _12815_/Y sky130_fd_sc_hd__o21ai_1
X_15534_ _15534_/A _15534_/B VGND VGND VPWR VPWR _15534_/Y sky130_fd_sc_hd__nand2_1
X_13795_ _13796_/A _13796_/B VGND VGND VPWR VPWR _13795_/X sky130_fd_sc_hd__and2_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12746_ _12697_/A _12697_/B _12697_/Y VGND VGND VPWR VPWR _12746_/X sky130_fd_sc_hd__a21o_1
XFILLER_42_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15465_ _15465_/A _15400_/X VGND VGND VPWR VPWR _15465_/X sky130_fd_sc_hd__or2b_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _12677_/A VGND VGND VPWR VPWR _12677_/Y sky130_fd_sc_hd__inv_2
X_15396_ _15396_/A _15396_/B VGND VGND VPWR VPWR _15471_/A sky130_fd_sc_hd__and2_1
X_14416_ _15030_/A _11742_/Y _11780_/Y _14415_/Y VGND VGND VPWR VPWR _14416_/X sky130_fd_sc_hd__o22a_1
X_11628_ _12413_/A _11627_/B _11627_/Y VGND VGND VPWR VPWR _11628_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14347_ _14381_/A _15952_/A VGND VGND VPWR VPWR _14347_/X sky130_fd_sc_hd__and2_1
XFILLER_7_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11559_ _11483_/X _11558_/X _11483_/X _11558_/X VGND VGND VPWR VPWR _11561_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14278_ _14179_/Y _14276_/Y _14277_/Y VGND VGND VPWR VPWR _14285_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16017_ _15939_/X _16017_/B VGND VGND VPWR VPWR _16017_/Y sky130_fd_sc_hd__nand2b_1
X_13229_ _13199_/X _13228_/Y _13199_/X _13228_/Y VGND VGND VPWR VPWR _13297_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _08770_/A _10132_/A VGND VGND VPWR VPWR _08770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09322_ _09322_/A VGND VGND VPWR VPWR _09327_/A sky130_fd_sc_hd__inv_2
XFILLER_40_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09253_ _08916_/A _10102_/B _08935_/X _08935_/A _08935_/B VGND VGND VPWR VPWR _09300_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09184_ _09184_/A VGND VGND VPWR VPWR _09184_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08968_ _08968_/A _08968_/B VGND VGND VPWR VPWR _08968_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08899_ _10014_/A _10128_/A _08803_/Y VGND VGND VPWR VPWR _08899_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10930_ _09322_/A _10928_/A _09327_/A _10928_/Y _11586_/A VGND VGND VPWR VPWR _12106_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_83_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12600_ _12595_/Y _12599_/A _12595_/A _12599_/Y _11708_/A VGND VGND VPWR VPWR _12618_/A
+ sky130_fd_sc_hd__o221a_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10861_ _10777_/X _10860_/Y _10777_/X _10860_/Y VGND VGND VPWR VPWR _10919_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10792_ _10791_/Y _10655_/X _10702_/Y VGND VGND VPWR VPWR _10792_/X sky130_fd_sc_hd__o21a_1
X_13580_ _12851_/A _13547_/B _13548_/Y _13579_/X VGND VGND VPWR VPWR _13580_/X sky130_fd_sc_hd__o22a_1
XFILLER_25_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ _13439_/A _11379_/B _11379_/Y VGND VGND VPWR VPWR _12532_/B sky130_fd_sc_hd__o21a_1
X_15250_ _15196_/A _15196_/B _15196_/Y VGND VGND VPWR VPWR _15250_/Y sky130_fd_sc_hd__o21ai_1
X_12462_ _15285_/A _12462_/B VGND VGND VPWR VPWR _12464_/B sky130_fd_sc_hd__or2_1
XFILLER_40_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14201_ _14201_/A _12628_/X VGND VGND VPWR VPWR _14201_/X sky130_fd_sc_hd__or2b_1
X_11413_ _11413_/A _11413_/B _12234_/B VGND VGND VPWR VPWR _12237_/A sky130_fd_sc_hd__or3_1
XFILLER_8_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15181_ _15181_/A _15181_/B VGND VGND VPWR VPWR _15181_/Y sky130_fd_sc_hd__nand2_1
X_12393_ _12393_/A _12456_/B VGND VGND VPWR VPWR _12393_/Y sky130_fd_sc_hd__nand2_1
X_14132_ _14132_/A VGND VGND VPWR VPWR _14132_/Y sky130_fd_sc_hd__inv_2
X_11344_ _13792_/A _11493_/B _11343_/Y VGND VGND VPWR VPWR _11344_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14063_ _14063_/A _14063_/B VGND VGND VPWR VPWR _14134_/B sky130_fd_sc_hd__or2_1
X_11275_ _11275_/A VGND VGND VPWR VPWR _12859_/A sky130_fd_sc_hd__buf_1
XFILLER_4_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13014_ _13014_/A VGND VGND VPWR VPWR _14496_/A sky130_fd_sc_hd__buf_1
X_10226_ _10226_/A VGND VGND VPWR VPWR _10226_/X sky130_fd_sc_hd__buf_1
XFILLER_121_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10157_ _10159_/A VGND VGND VPWR VPWR _10243_/B sky130_fd_sc_hd__buf_1
X_14965_ _15563_/A _14982_/B _14964_/Y VGND VGND VPWR VPWR _14965_/Y sky130_fd_sc_hd__o21ai_1
X_10088_ _10037_/X _10086_/X _11523_/B VGND VGND VPWR VPWR _10088_/X sky130_fd_sc_hd__o21a_1
X_13916_ _15406_/A _13947_/B VGND VGND VPWR VPWR _13916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14896_ _14809_/A _14809_/B _14809_/Y VGND VGND VPWR VPWR _14896_/X sky130_fd_sc_hd__a21o_1
XFILLER_90_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13847_ _14622_/A _13847_/B VGND VGND VPWR VPWR _13847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13778_ _15116_/A _13778_/B VGND VGND VPWR VPWR _13778_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15517_ _15467_/A _15467_/B _15467_/Y VGND VGND VPWR VPWR _15517_/Y sky130_fd_sc_hd__o21ai_1
X_12729_ _12719_/X _12728_/X _12719_/X _12728_/X VGND VGND VPWR VPWR _12784_/B sky130_fd_sc_hd__a2bb2o_1
X_15448_ _15411_/X _15447_/X _15411_/X _15447_/X VGND VGND VPWR VPWR _15449_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15379_ _15338_/X _15378_/X _15338_/X _15378_/X VGND VGND VPWR VPWR _15406_/B sky130_fd_sc_hd__a2bb2o_1
X_09940_ _11595_/A VGND VGND VPWR VPWR _09941_/A sky130_fd_sc_hd__inv_2
XFILLER_98_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09871_ _09449_/Y _09870_/X _09476_/X VGND VGND VPWR VPWR _09871_/X sky130_fd_sc_hd__o21a_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _08822_/A VGND VGND VPWR VPWR _08823_/A sky130_fd_sc_hd__inv_2
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _09478_/A _10134_/A _08752_/X VGND VGND VPWR VPWR _08753_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_81_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08684_ _09549_/A _08609_/A _08611_/Y _08683_/X VGND VGND VPWR VPWR _08684_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09305_ _10245_/A _09306_/B VGND VGND VPWR VPWR _09305_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09236_ _08721_/B _09799_/A _09231_/Y _09628_/A VGND VGND VPWR VPWR _09237_/A sky130_fd_sc_hd__o22a_1
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09167_ _10008_/B _09167_/B VGND VGND VPWR VPWR _09167_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09098_ _09409_/A VGND VGND VPWR VPWR _09714_/A sky130_fd_sc_hd__inv_2
XFILLER_119_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11060_ _12234_/A VGND VGND VPWR VPWR _11795_/A sky130_fd_sc_hd__inv_2
XFILLER_1_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10011_ _10011_/A _10011_/B VGND VGND VPWR VPWR _10041_/B sky130_fd_sc_hd__nor2_1
XFILLER_130_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14750_ _14676_/A _14676_/B _14669_/X _14676_/Y VGND VGND VPWR VPWR _14750_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11962_ _13004_/A _11893_/B _11893_/Y VGND VGND VPWR VPWR _11962_/Y sky130_fd_sc_hd__o21ai_1
X_13701_ _13726_/A _13699_/X _13700_/X VGND VGND VPWR VPWR _13701_/X sky130_fd_sc_hd__o21a_1
XFILLER_57_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10913_ _10901_/Y _10911_/X _10912_/Y VGND VGND VPWR VPWR _10913_/X sky130_fd_sc_hd__o21a_1
X_14681_ _14681_/A _14680_/X VGND VGND VPWR VPWR _14681_/X sky130_fd_sc_hd__or2b_1
X_11893_ _13004_/A _11893_/B VGND VGND VPWR VPWR _11893_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16420_ _16437_/B _16429_/B VGND VGND VPWR VPWR _16420_/X sky130_fd_sc_hd__or2_1
XFILLER_71_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10844_ _10939_/A _10843_/Y _10939_/A _10843_/Y VGND VGND VPWR VPWR _10845_/B sky130_fd_sc_hd__a2bb2o_1
X_13632_ _13632_/A VGND VGND VPWR VPWR _15128_/A sky130_fd_sc_hd__buf_1
XFILLER_44_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16351_ _16334_/A _16334_/B _16334_/Y VGND VGND VPWR VPWR _16351_/Y sky130_fd_sc_hd__o21ai_1
X_13563_ _13563_/A _13563_/B VGND VGND VPWR VPWR _13564_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12514_ _14131_/A VGND VGND VPWR VPWR _13443_/A sky130_fd_sc_hd__buf_1
X_15302_ _15347_/A _15347_/B VGND VGND VPWR VPWR _15366_/A sky130_fd_sc_hd__and2_1
X_10775_ _13083_/A _10741_/B _10741_/Y _10774_/X VGND VGND VPWR VPWR _10775_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16282_ _16270_/A _16336_/A _16270_/Y VGND VGND VPWR VPWR _16282_/Y sky130_fd_sc_hd__o21ai_1
X_13494_ _13494_/A _13494_/B VGND VGND VPWR VPWR _13494_/X sky130_fd_sc_hd__and2_1
XFILLER_13_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12445_ _12445_/A VGND VGND VPWR VPWR _15285_/A sky130_fd_sc_hd__clkbuf_2
X_15233_ _15228_/X _15232_/Y _15228_/X _15232_/Y VGND VGND VPWR VPWR _15234_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15164_ _12431_/A _15163_/B _15163_/Y VGND VGND VPWR VPWR _15164_/X sky130_fd_sc_hd__a21o_1
X_12376_ _12376_/A _12376_/B VGND VGND VPWR VPWR _12376_/X sky130_fd_sc_hd__or2_1
X_14115_ _14078_/Y _14112_/X _14880_/A _14114_/Y VGND VGND VPWR VPWR _14115_/X sky130_fd_sc_hd__o22a_1
X_11327_ _11521_/A _11521_/B _11326_/Y VGND VGND VPWR VPWR _11328_/A sky130_fd_sc_hd__o21ai_2
XFILLER_4_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15095_ _15066_/A _15066_/B _15066_/Y _15094_/X VGND VGND VPWR VPWR _15095_/X sky130_fd_sc_hd__a2bb2o_1
X_14046_ _14046_/A VGND VGND VPWR VPWR _14046_/X sky130_fd_sc_hd__buf_1
X_11258_ _14027_/A _11219_/B _11219_/Y _11257_/X VGND VGND VPWR VPWR _11258_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10209_ _10906_/A _10215_/A VGND VGND VPWR VPWR _10210_/A sky130_fd_sc_hd__or2_1
X_11189_ _09426_/A _09136_/B _09136_/Y VGND VGND VPWR VPWR _11190_/A sky130_fd_sc_hd__o21ai_1
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15997_ _15969_/Y _15996_/X _15969_/Y _15996_/X VGND VGND VPWR VPWR _16053_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14948_ _14948_/A _14948_/B VGND VGND VPWR VPWR _14948_/X sky130_fd_sc_hd__or2_1
X_14879_ _15544_/A _14920_/B VGND VGND VPWR VPWR _14879_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09021_ _08580_/X _08893_/X _09021_/S VGND VGND VPWR VPWR _09553_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09923_ _09923_/A _09923_/B VGND VGND VPWR VPWR _11300_/A sky130_fd_sc_hd__nor2_1
X_09854_ _09855_/A _09854_/B VGND VGND VPWR VPWR _09854_/Y sky130_fd_sc_hd__nor2_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08805_ _08794_/A _09467_/B _08714_/Y VGND VGND VPWR VPWR _08806_/A sky130_fd_sc_hd__a21oi_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09785_ _09785_/A _09785_/B VGND VGND VPWR VPWR _09785_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08736_ _08736_/A VGND VGND VPWR VPWR _08736_/Y sky130_fd_sc_hd__inv_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08667_ _08667_/A VGND VGND VPWR VPWR _08667_/Y sky130_fd_sc_hd__inv_2
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08598_ _08598_/A VGND VGND VPWR VPWR _08598_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10560_ _10968_/A _11207_/A VGND VGND VPWR VPWR _10561_/A sky130_fd_sc_hd__or2_1
X_10491_ _10489_/Y _10490_/Y _10490_/A _09847_/B _09941_/A VGND VGND VPWR VPWR _12930_/A
+ sky130_fd_sc_hd__o221a_2
X_09219_ _09549_/A _09696_/A VGND VGND VPWR VPWR _09220_/A sky130_fd_sc_hd__or2_1
XFILLER_108_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12230_ _12230_/A _12139_/X VGND VGND VPWR VPWR _12230_/X sky130_fd_sc_hd__or2b_1
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12161_ _12160_/Y _12069_/X _12103_/Y VGND VGND VPWR VPWR _12161_/X sky130_fd_sc_hd__o21a_1
X_12092_ _12780_/A _12170_/A VGND VGND VPWR VPWR _12092_/Y sky130_fd_sc_hd__nor2_1
X_11112_ _09661_/X _11111_/X _09661_/X _11111_/X VGND VGND VPWR VPWR _11113_/B sky130_fd_sc_hd__a2bb2oi_1
X_15920_ _15901_/X _15919_/Y _15901_/X _15919_/Y VGND VGND VPWR VPWR _15964_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11043_ _12843_/A VGND VGND VPWR VPWR _15078_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15851_ _14283_/A _15850_/X _12638_/X VGND VGND VPWR VPWR _15851_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14802_ _14802_/A _14802_/B VGND VGND VPWR VPWR _14802_/X sky130_fd_sc_hd__and2_1
XFILLER_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15782_ _14363_/A _15777_/A _14375_/A VGND VGND VPWR VPWR _16028_/B sky130_fd_sc_hd__a21bo_1
X_12994_ _14462_/A _12930_/B _12930_/Y VGND VGND VPWR VPWR _12994_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14733_ _14792_/A _14731_/X _14732_/X VGND VGND VPWR VPWR _14733_/X sky130_fd_sc_hd__o21a_1
X_11945_ _11976_/A _11976_/B VGND VGND VPWR VPWR _11945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14664_ _14664_/A _14664_/B VGND VGND VPWR VPWR _14664_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16403_ _16393_/Y _16401_/X _16349_/X _16402_/X VGND VGND VPWR VPWR _16404_/B sky130_fd_sc_hd__o31a_1
X_13615_ _13615_/A VGND VGND VPWR VPWR _13615_/Y sky130_fd_sc_hd__inv_2
X_11876_ _11907_/A _11907_/B VGND VGND VPWR VPWR _11876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14595_ _12093_/Y _14594_/X _12093_/Y _14594_/X VGND VGND VPWR VPWR _14596_/B sky130_fd_sc_hd__o2bb2a_1
X_10827_ _10815_/X _10826_/Y _10815_/X _10826_/Y VGND VGND VPWR VPWR _10964_/A sky130_fd_sc_hd__o2bb2a_1
X_16334_ _16334_/A _16334_/B VGND VGND VPWR VPWR _16334_/Y sky130_fd_sc_hd__nand2_1
X_10758_ _10763_/A _10758_/B VGND VGND VPWR VPWR _13752_/A sky130_fd_sc_hd__or2_1
X_13546_ _13536_/X _13545_/Y _13536_/X _13545_/Y VGND VGND VPWR VPWR _13547_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16265_ _16178_/Y _16263_/X _16264_/Y VGND VGND VPWR VPWR _16265_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13477_ _14308_/A _13477_/B VGND VGND VPWR VPWR _15982_/A sky130_fd_sc_hd__or2_1
XFILLER_9_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15216_ _15216_/A _15216_/B VGND VGND VPWR VPWR _15216_/X sky130_fd_sc_hd__or2_1
X_12428_ _12428_/A VGND VGND VPWR VPWR _12429_/A sky130_fd_sc_hd__inv_2
X_10689_ _10689_/A VGND VGND VPWR VPWR _10689_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_126_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16196_ _16196_/A VGND VGND VPWR VPWR _16196_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12359_ _12295_/X _12250_/X _12297_/B VGND VGND VPWR VPWR _12359_/X sky130_fd_sc_hd__o21a_1
X_15147_ _15146_/A _15146_/B _10522_/Y _15146_/Y VGND VGND VPWR VPWR _15147_/X sky130_fd_sc_hd__a2bb2o_1
X_15078_ _15078_/A _15078_/B VGND VGND VPWR VPWR _15078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14029_ _15404_/A _13945_/B _13945_/Y VGND VGND VPWR VPWR _14029_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09570_ _09482_/A _09482_/B _09482_/Y VGND VGND VPWR VPWR _09570_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08521_ _08697_/A _08521_/B VGND VGND VPWR VPWR _09862_/A sky130_fd_sc_hd__or2_1
XFILLER_35_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08452_ _08543_/B _08446_/Y _09331_/A VGND VGND VPWR VPWR _08453_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08383_ _08642_/A VGND VGND VPWR VPWR _09228_/A sky130_fd_sc_hd__buf_1
XFILLER_51_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09004_ _12302_/A VGND VGND VPWR VPWR _14137_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09906_ _10657_/A _10656_/A VGND VGND VPWR VPWR _09907_/B sky130_fd_sc_hd__or2_1
XFILLER_116_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09837_ _09832_/A _09832_/B _09833_/Y _09836_/Y VGND VGND VPWR VPWR _09838_/B sky130_fd_sc_hd__o22a_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09768_ _10052_/A VGND VGND VPWR VPWR _10077_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08719_ _08944_/A _08719_/B VGND VGND VPWR VPWR _08719_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11730_ _11787_/A _11722_/B _11722_/Y _11787_/B VGND VGND VPWR VPWR _11731_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09699_ _09698_/A _09698_/B _09730_/A VGND VGND VPWR VPWR _09700_/A sky130_fd_sc_hd__a21bo_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _12789_/A _11661_/B VGND VGND VPWR VPWR _11661_/X sky130_fd_sc_hd__or2_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14380_ _14353_/X _14378_/X _15644_/B VGND VGND VPWR VPWR _14380_/X sky130_fd_sc_hd__o21a_1
X_13400_ _14090_/A VGND VGND VPWR VPWR _14908_/A sky130_fd_sc_hd__buf_1
X_10612_ _11888_/A VGND VGND VPWR VPWR _11895_/A sky130_fd_sc_hd__buf_1
X_11592_ _09789_/X _11591_/Y _09789_/X _11591_/Y VGND VGND VPWR VPWR _11593_/B sky130_fd_sc_hd__a2bb2oi_1
X_13331_ _13331_/A _13331_/B VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__and2_1
X_10543_ _10543_/A _10543_/B VGND VGND VPWR VPWR _10543_/Y sky130_fd_sc_hd__nand2_1
X_16050_ _15968_/X _16049_/Y _15968_/X _16049_/Y VGND VGND VPWR VPWR _16050_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13262_ _13824_/A _13186_/B _13186_/Y VGND VGND VPWR VPWR _13262_/Y sky130_fd_sc_hd__o21ai_1
X_15001_ _11766_/X _15000_/X _11768_/B VGND VGND VPWR VPWR _15001_/X sky130_fd_sc_hd__o21a_1
X_10474_ _10554_/A _11855_/A VGND VGND VPWR VPWR _10474_/Y sky130_fd_sc_hd__nor2_1
X_12213_ _12150_/X _12212_/X _12150_/X _12212_/X VGND VGND VPWR VPWR _12214_/B sky130_fd_sc_hd__a2bb2o_1
X_13193_ _13165_/Y _13191_/X _13192_/Y VGND VGND VPWR VPWR _13193_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12144_ _12224_/A _12142_/X _12143_/X VGND VGND VPWR VPWR _12144_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12075_ _13583_/A _12075_/B VGND VGND VPWR VPWR _12075_/X sky130_fd_sc_hd__and2_1
XFILLER_1_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15903_ _15859_/Y _15901_/X _15902_/Y VGND VGND VPWR VPWR _15906_/B sky130_fd_sc_hd__o21a_1
XFILLER_110_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11026_ _15069_/A VGND VGND VPWR VPWR _13909_/A sky130_fd_sc_hd__buf_1
XFILLER_77_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15834_ _15706_/X _15834_/B VGND VGND VPWR VPWR _15834_/X sky130_fd_sc_hd__and2b_1
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15765_ _14907_/X _15764_/X _14907_/X _15764_/X VGND VGND VPWR VPWR _15766_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12977_ _14476_/A _12938_/B _12938_/Y VGND VGND VPWR VPWR _12977_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15696_ _16055_/A _15696_/B VGND VGND VPWR VPWR _15696_/Y sky130_fd_sc_hd__nand2_1
X_14716_ _14644_/Y _14715_/X _14644_/Y _14715_/X VGND VGND VPWR VPWR _14717_/B sky130_fd_sc_hd__a2bb2o_1
X_11928_ _11928_/A _11928_/B VGND VGND VPWR VPWR _11929_/B sky130_fd_sc_hd__or2_1
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14647_ _15333_/A _14647_/B VGND VGND VPWR VPWR _14647_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11859_ _11859_/A VGND VGND VPWR VPWR _11923_/B sky130_fd_sc_hd__inv_2
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14578_ _14558_/Y _14576_/X _14577_/Y VGND VGND VPWR VPWR _14578_/X sky130_fd_sc_hd__o21a_1
X_16317_ _16312_/Y _16315_/Y _16316_/Y VGND VGND VPWR VPWR _16317_/X sky130_fd_sc_hd__o21a_1
X_13529_ _13529_/A _13529_/B VGND VGND VPWR VPWR _13529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16248_ _16457_/S _16248_/B VGND VGND VPWR VPWR _16248_/Y sky130_fd_sc_hd__nor2_1
X_16179_ _16076_/X _16179_/B VGND VGND VPWR VPWR _16179_/X sky130_fd_sc_hd__and2b_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09622_ _09502_/A _09502_/B _09502_/Y VGND VGND VPWR VPWR _09622_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09553_ _09553_/A _09553_/B VGND VGND VPWR VPWR _09601_/B sky130_fd_sc_hd__and2_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08504_ _09448_/B VGND VGND VPWR VPWR _09561_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09484_ _09484_/A _09484_/B VGND VGND VPWR VPWR _09484_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08435_ _08434_/A _08328_/Y _08434_/Y _08328_/A _08441_/A VGND VGND VPWR VPWR _10012_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08366_ _08366_/A VGND VGND VPWR VPWR _08366_/Y sky130_fd_sc_hd__inv_2
X_08297_ input24/X input8/X input24/X input8/X VGND VGND VPWR VPWR _08298_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_133_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10190_ _10240_/B _10147_/B _10147_/Y _10189_/X VGND VGND VPWR VPWR _10190_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13880_ _13862_/X _13879_/Y _13862_/X _13879_/Y VGND VGND VPWR VPWR _13882_/B sky130_fd_sc_hd__a2bb2o_1
X_12900_ _14464_/A _12932_/B VGND VGND VPWR VPWR _12900_/Y sky130_fd_sc_hd__nor2_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _12830_/A _12830_/B _12830_/Y VGND VGND VPWR VPWR _12831_/X sky130_fd_sc_hd__a21o_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _15550_/A _15550_/B VGND VGND VPWR VPWR _15690_/B sky130_fd_sc_hd__or2_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12762_ _10342_/X _10424_/B _10342_/X _10424_/B VGND VGND VPWR VPWR _12833_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _14790_/A _15452_/B _15452_/X _15480_/X VGND VGND VPWR VPWR _15481_/X sky130_fd_sc_hd__o22a_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14458_/A _14458_/B _14458_/Y VGND VGND VPWR VPWR _14501_/X sky130_fd_sc_hd__o21a_1
X_11713_ _11713_/A VGND VGND VPWR VPWR _11774_/A sky130_fd_sc_hd__clkinvlp_2
X_12693_ _12693_/A _12693_/B VGND VGND VPWR VPWR _12693_/Y sky130_fd_sc_hd__nor2_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _12141_/A _14426_/B _14426_/X _14431_/X VGND VGND VPWR VPWR _14432_/X sky130_fd_sc_hd__o22a_1
X_11644_ _12454_/A _11644_/B VGND VGND VPWR VPWR _11644_/X sky130_fd_sc_hd__or2_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 wbs_dat_i[3] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__buf_4
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14363_ _14363_/A _15777_/A VGND VGND VPWR VPWR _14375_/A sky130_fd_sc_hd__or2_1
X_16102_ _16036_/A _16036_/B _16036_/Y VGND VGND VPWR VPWR _16102_/Y sky130_fd_sc_hd__o21ai_1
X_11575_ _14065_/A VGND VGND VPWR VPWR _15437_/A sky130_fd_sc_hd__buf_1
Xinput16 wbs_adr_i[8] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_2
XFILLER_116_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14294_ _14172_/X _14294_/B VGND VGND VPWR VPWR _14294_/Y sky130_fd_sc_hd__nand2b_1
X_13314_ _14771_/A _13303_/B _13303_/Y VGND VGND VPWR VPWR _13314_/Y sky130_fd_sc_hd__o21ai_1
X_10526_ _10513_/Y _10524_/X _10525_/Y VGND VGND VPWR VPWR _10526_/X sky130_fd_sc_hd__o21a_1
X_16033_ _16022_/Y _16031_/X _16032_/Y VGND VGND VPWR VPWR _16033_/X sky130_fd_sc_hd__o21a_1
X_13245_ _14732_/A _13288_/B VGND VGND VPWR VPWR _13245_/Y sky130_fd_sc_hd__nor2_1
X_10457_ _10968_/A _11214_/A VGND VGND VPWR VPWR _10458_/A sky130_fd_sc_hd__or2_1
XFILLER_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13176_ _14563_/A _13103_/B _13103_/Y VGND VGND VPWR VPWR _13176_/Y sky130_fd_sc_hd__o21ai_1
X_10388_ _10450_/A _12699_/A _10387_/Y VGND VGND VPWR VPWR _10388_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12127_ _13921_/A _12143_/B VGND VGND VPWR VPWR _12224_/A sky130_fd_sc_hd__and2_1
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12058_ _12032_/Y _12056_/X _12057_/Y VGND VGND VPWR VPWR _12058_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11009_ _11009_/A VGND VGND VPWR VPWR _13583_/A sky130_fd_sc_hd__buf_1
XFILLER_38_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15817_ _15817_/A _15817_/B VGND VGND VPWR VPWR _15817_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15748_ _15676_/X _15747_/Y _15676_/X _15747_/Y VGND VGND VPWR VPWR _15809_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15679_ _15679_/A _15679_/B VGND VGND VPWR VPWR _15679_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08984_ _08984_/A _08984_/B VGND VGND VPWR VPWR _11462_/B sky130_fd_sc_hd__or2_1
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09605_ _09510_/X _09604_/X _09510_/X _09604_/X VGND VGND VPWR VPWR _09980_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09536_ _09549_/A _09549_/B VGND VGND VPWR VPWR _09613_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09467_ _10014_/A _09467_/B VGND VGND VPWR VPWR _09467_/X sky130_fd_sc_hd__or2_1
XFILLER_24_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08418_ _08418_/A VGND VGND VPWR VPWR _08418_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09398_ _15060_/A VGND VGND VPWR VPWR _13897_/A sky130_fd_sc_hd__buf_1
X_08349_ _08349_/A VGND VGND VPWR VPWR _08349_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11360_ _08979_/X _11359_/X _08979_/X _11359_/X VGND VGND VPWR VPWR _11361_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_125_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10311_ _10309_/A _10309_/B _10310_/A _10309_/Y _10310_/Y VGND VGND VPWR VPWR _10367_/A
+ sky130_fd_sc_hd__o32a_1
X_13030_ _13055_/A _13028_/X _13029_/X VGND VGND VPWR VPWR _13030_/X sky130_fd_sc_hd__o21a_1
X_11291_ _11291_/A VGND VGND VPWR VPWR _11291_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10242_ _10242_/A _10242_/B VGND VGND VPWR VPWR _10242_/X sky130_fd_sc_hd__or2_1
XFILLER_121_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10173_ _10173_/A _10173_/B VGND VGND VPWR VPWR _10173_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14981_ _14980_/Y _14945_/X _14942_/Y VGND VGND VPWR VPWR _14981_/X sky130_fd_sc_hd__o21a_1
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13932_ _14429_/A VGND VGND VPWR VPWR _15396_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13863_ _13863_/A VGND VGND VPWR VPWR _13863_/Y sky130_fd_sc_hd__inv_2
X_15602_ _15602_/A VGND VGND VPWR VPWR _15602_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_74_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13794_ _13776_/X _13793_/Y _13776_/X _13793_/Y VGND VGND VPWR VPWR _13796_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12814_ _12847_/A _12847_/B VGND VGND VPWR VPWR _12814_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15533_ _15478_/X _15532_/Y _15478_/X _15532_/Y VGND VGND VPWR VPWR _15616_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _12774_/A _12774_/B VGND VGND VPWR VPWR _12745_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15464_ _15464_/A _15464_/B VGND VGND VPWR VPWR _15464_/Y sky130_fd_sc_hd__nand2_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _11521_/Y _12675_/Y _11326_/Y VGND VGND VPWR VPWR _12677_/A sky130_fd_sc_hd__o21ai_2
X_15395_ _15396_/A _15396_/B VGND VGND VPWR VPWR _15395_/X sky130_fd_sc_hd__or2_1
X_14415_ _14415_/A VGND VGND VPWR VPWR _14415_/Y sky130_fd_sc_hd__inv_2
X_11627_ _12413_/A _11627_/B VGND VGND VPWR VPWR _11627_/Y sky130_fd_sc_hd__nor2_1
X_14346_ _14352_/A _14346_/B VGND VGND VPWR VPWR _15952_/A sky130_fd_sc_hd__or2_1
X_11558_ _11558_/A _11557_/X VGND VGND VPWR VPWR _11558_/X sky130_fd_sc_hd__or2b_1
XFILLER_116_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10509_ _13608_/A VGND VGND VPWR VPWR _11838_/A sky130_fd_sc_hd__inv_2
XFILLER_7_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16016_ _16036_/A _16036_/B VGND VGND VPWR VPWR _16016_/Y sky130_fd_sc_hd__nor2_1
X_14277_ _14277_/A _14277_/B VGND VGND VPWR VPWR _14277_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11489_ _09997_/A _09666_/B _09666_/Y VGND VGND VPWR VPWR _11489_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13228_ _13200_/A _13200_/B _13200_/Y VGND VGND VPWR VPWR _13228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13159_ _13196_/A _13196_/B VGND VGND VPWR VPWR _13159_/Y sky130_fd_sc_hd__nor2_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09321_ _09318_/X _09320_/X _09318_/X _09320_/X VGND VGND VPWR VPWR _09322_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09252_ _09458_/A _09252_/B VGND VGND VPWR VPWR _10061_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09183_ _09525_/B _09156_/B _09156_/X VGND VGND VPWR VPWR _09184_/A sky130_fd_sc_hd__a21bo_1
XFILLER_108_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08967_ _08682_/X _08966_/X _08682_/X _08966_/X VGND VGND VPWR VPWR _11395_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08898_ _08685_/X _08897_/X _08685_/X _08897_/X VGND VGND VPWR VPWR _08974_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10860_ _11976_/A _10716_/B _10716_/Y VGND VGND VPWR VPWR _10860_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09519_ _09518_/A _09518_/B _09563_/A _09518_/X VGND VGND VPWR VPWR _09519_/Y sky130_fd_sc_hd__o22ai_1
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10791_ _13636_/A _10791_/B VGND VGND VPWR VPWR _10791_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _14119_/A VGND VGND VPWR VPWR _13439_/A sky130_fd_sc_hd__buf_1
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12461_ _12460_/Y _12363_/Y _12396_/Y VGND VGND VPWR VPWR _12461_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14200_ _14206_/A _14200_/B VGND VGND VPWR VPWR _15866_/A sky130_fd_sc_hd__or2_1
X_11412_ _12322_/A VGND VGND VPWR VPWR _13405_/A sky130_fd_sc_hd__inv_2
X_15180_ _15157_/X _15179_/Y _15157_/X _15179_/Y VGND VGND VPWR VPWR _15181_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14131_ _14131_/A VGND VGND VPWR VPWR _14868_/A sky130_fd_sc_hd__inv_2
X_12392_ _12368_/X _12391_/Y _12368_/X _12391_/Y VGND VGND VPWR VPWR _12456_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11343_ _12364_/A _11493_/B VGND VGND VPWR VPWR _11343_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14062_ _14011_/X _14060_/X _14128_/B VGND VGND VPWR VPWR _14062_/X sky130_fd_sc_hd__o21a_1
X_11274_ _13785_/A VGND VGND VPWR VPWR _11275_/A sky130_fd_sc_hd__buf_1
XFILLER_121_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13013_ _13003_/Y _13011_/X _13012_/Y VGND VGND VPWR VPWR _13013_/X sky130_fd_sc_hd__o21a_1
X_10225_ _10224_/A _10224_/B _10309_/A VGND VGND VPWR VPWR _10226_/A sky130_fd_sc_hd__o21bai_1
XFILLER_121_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10156_ _10115_/A _10115_/B _10116_/A VGND VGND VPWR VPWR _10159_/A sky130_fd_sc_hd__a21bo_1
X_14964_ _15563_/A _14982_/B VGND VGND VPWR VPWR _14964_/Y sky130_fd_sc_hd__nand2_1
X_10087_ _10087_/A _10087_/B VGND VGND VPWR VPWR _11523_/B sky130_fd_sc_hd__or2_1
X_13915_ _13846_/X _13914_/Y _13846_/X _13914_/Y VGND VGND VPWR VPWR _13947_/B sky130_fd_sc_hd__a2bb2o_1
X_14895_ _15524_/A _14910_/B VGND VGND VPWR VPWR _14895_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13846_ _13820_/Y _13844_/X _13845_/Y VGND VGND VPWR VPWR _13846_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13777_ _13777_/A VGND VGND VPWR VPWR _13777_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10989_ _10965_/X _10988_/X _10965_/X _10988_/X VGND VGND VPWR VPWR _11130_/B sky130_fd_sc_hd__a2bb2o_1
X_15516_ _15519_/A _15519_/B VGND VGND VPWR VPWR _15639_/A sky130_fd_sc_hd__and2_1
XFILLER_43_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12728_ _12685_/A _12685_/B _12685_/Y VGND VGND VPWR VPWR _12728_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15447_ _15447_/A _15412_/X VGND VGND VPWR VPWR _15447_/X sky130_fd_sc_hd__or2b_1
X_12659_ _10224_/A _10224_/B _12658_/Y VGND VGND VPWR VPWR _12659_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15378_ _15378_/A _15339_/X VGND VGND VPWR VPWR _15378_/X sky130_fd_sc_hd__or2b_1
X_14329_ _14387_/A _15958_/A VGND VGND VPWR VPWR _14329_/X sky130_fd_sc_hd__and2_1
XFILLER_116_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09870_ _09450_/Y _09869_/X _09474_/X VGND VGND VPWR VPWR _09870_/X sky130_fd_sc_hd__o21a_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08821_ _09221_/A _09456_/B _08716_/X VGND VGND VPWR VPWR _08822_/A sky130_fd_sc_hd__o21ai_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _10008_/A _10134_/A VGND VGND VPWR VPWR _08752_/X sky130_fd_sc_hd__or2_1
XFILLER_66_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08683_ _09547_/A _08622_/A _08624_/Y _08682_/X VGND VGND VPWR VPWR _08683_/X sky130_fd_sc_hd__o22a_1
XFILLER_81_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09304_ _10402_/A _09302_/Y _09303_/Y VGND VGND VPWR VPWR _09306_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09235_ _09629_/A VGND VGND VPWR VPWR _09628_/A sky130_fd_sc_hd__inv_2
X_09166_ _10009_/B _09166_/B VGND VGND VPWR VPWR _09167_/B sky130_fd_sc_hd__or2_1
XFILLER_134_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09097_ _09070_/A _09070_/B _09071_/B VGND VGND VPWR VPWR _09409_/A sky130_fd_sc_hd__a21bo_1
XFILLER_122_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10010_ _10010_/A _10010_/B VGND VGND VPWR VPWR _10038_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09999_ _09999_/A _09999_/B VGND VGND VPWR VPWR _10000_/A sky130_fd_sc_hd__nand2_1
X_11961_ _11961_/A VGND VGND VPWR VPWR _11961_/X sky130_fd_sc_hd__buf_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10912_ _13828_/A _10912_/B VGND VGND VPWR VPWR _10912_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13700_ _13700_/A _13700_/B VGND VGND VPWR VPWR _13700_/X sky130_fd_sc_hd__or2_1
XFILLER_57_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11892_ _11892_/A _11893_/B VGND VGND VPWR VPWR _11892_/Y sky130_fd_sc_hd__nor2_1
X_14680_ _15184_/A _14680_/B VGND VGND VPWR VPWR _14680_/X sky130_fd_sc_hd__or2_1
XFILLER_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10843_ _13700_/A _10938_/B _10842_/Y VGND VGND VPWR VPWR _10843_/Y sky130_fd_sc_hd__o21ai_1
X_13631_ _13631_/A VGND VGND VPWR VPWR _13631_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16350_ _08230_/X _16468_/Q _08233_/X _16349_/X _16343_/X VGND VGND VPWR VPWR _16468_/D
+ sky130_fd_sc_hd__o221a_2
X_10774_ _13088_/A _10749_/B _10749_/Y _10773_/X VGND VGND VPWR VPWR _10774_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13562_ _13532_/X _13561_/Y _13532_/X _13561_/Y VGND VGND VPWR VPWR _13563_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16281_ _16338_/A _16338_/B VGND VGND VPWR VPWR _16281_/Y sky130_fd_sc_hd__nor2_1
X_12513_ _12638_/A _12638_/B VGND VGND VPWR VPWR _14283_/A sky130_fd_sc_hd__and2_1
X_15301_ _15280_/X _15300_/Y _15280_/X _15300_/Y VGND VGND VPWR VPWR _15347_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13493_ _11620_/Y _13492_/X _11620_/Y _13492_/X VGND VGND VPWR VPWR _13494_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15232_ _15178_/A _15178_/B _15178_/Y VGND VGND VPWR VPWR _15232_/Y sky130_fd_sc_hd__o21ai_1
X_12444_ _13462_/A _12441_/B _12441_/X _12443_/X VGND VGND VPWR VPWR _12444_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12375_ _12437_/A VGND VGND VPWR VPWR _12786_/A sky130_fd_sc_hd__buf_1
X_15163_ _15163_/A _15163_/B VGND VGND VPWR VPWR _15163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14114_ _14114_/A VGND VGND VPWR VPWR _14114_/Y sky130_fd_sc_hd__inv_2
X_15094_ _15069_/A _15069_/B _15069_/Y _15093_/X VGND VGND VPWR VPWR _15094_/X sky130_fd_sc_hd__a2bb2o_1
X_11326_ _11521_/A _11521_/B VGND VGND VPWR VPWR _11326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14045_ _13936_/X _14044_/X _13936_/A _14044_/X VGND VGND VPWR VPWR _14047_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11257_ _14031_/A _11225_/B _11225_/Y _11256_/X VGND VGND VPWR VPWR _11257_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11188_ _14059_/A _11188_/B VGND VGND VPWR VPWR _11188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10208_ _10287_/A VGND VGND VPWR VPWR _10906_/A sky130_fd_sc_hd__inv_1
XFILLER_95_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10139_ _10139_/A _10139_/B VGND VGND VPWR VPWR _10139_/Y sky130_fd_sc_hd__nor2_1
X_15996_ _15970_/A _15970_/B _15970_/Y VGND VGND VPWR VPWR _15996_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14947_ _14948_/A _14948_/B VGND VGND VPWR VPWR _14949_/A sky130_fd_sc_hd__and2_1
XFILLER_63_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14878_ _14823_/X _14877_/X _14823_/X _14877_/X VGND VGND VPWR VPWR _14920_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13829_ _13756_/A _13756_/B _13756_/Y VGND VGND VPWR VPWR _13829_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09020_ _09470_/A _08567_/X _09020_/S VGND VGND VPWR VPWR _09555_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09922_ _09923_/A _09923_/B VGND VGND VPWR VPWR _11300_/B sky130_fd_sc_hd__and2_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09853_ _09853_/A _09853_/B VGND VGND VPWR VPWR _09854_/B sky130_fd_sc_hd__and2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08804_ _09249_/A VGND VGND VPWR VPWR _09494_/A sky130_fd_sc_hd__buf_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _09785_/A _09785_/B VGND VGND VPWR VPWR _09784_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08735_ _08712_/Y _08733_/Y _08734_/X VGND VGND VPWR VPWR _08736_/A sky130_fd_sc_hd__o21ai_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08666_ _08666_/A1 _08398_/A _09232_/A _08398_/Y VGND VGND VPWR VPWR _08667_/A sky130_fd_sc_hd__o22a_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08597_ _08597_/A _10114_/B VGND VGND VPWR VPWR _08598_/A sky130_fd_sc_hd__or2_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10490_ _10490_/A _10490_/B VGND VGND VPWR VPWR _10490_/Y sky130_fd_sc_hd__nor2_1
X_09218_ _09803_/A VGND VGND VPWR VPWR _09696_/A sky130_fd_sc_hd__inv_2
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09149_ _09518_/A _09148_/X _08521_/B VGND VGND VPWR VPWR _09150_/S sky130_fd_sc_hd__o21ba_1
X_12160_ _13053_/A _12160_/B VGND VGND VPWR VPWR _12160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11111_ _09993_/A _09662_/B _09662_/Y VGND VGND VPWR VPWR _11111_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12091_ _12174_/B _12090_/X _12174_/B _12090_/X VGND VGND VPWR VPWR _12170_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11042_ _13563_/A VGND VGND VPWR VPWR _12843_/A sky130_fd_sc_hd__buf_1
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15850_ _14177_/A _15849_/X _12636_/X VGND VGND VPWR VPWR _15850_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14801_ _14727_/X _14800_/X _14727_/X _14800_/X VGND VGND VPWR VPWR _14802_/B sky130_fd_sc_hd__a2bb2o_1
X_15781_ _15781_/A _15781_/B VGND VGND VPWR VPWR _15784_/A sky130_fd_sc_hd__nor2_1
XFILLER_92_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12993_ _13672_/A VGND VGND VPWR VPWR _14492_/A sky130_fd_sc_hd__buf_1
XFILLER_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14732_ _14732_/A _14732_/B VGND VGND VPWR VPWR _14732_/X sky130_fd_sc_hd__or2_1
X_11944_ _11909_/A _11943_/Y _11909_/A _11943_/Y VGND VGND VPWR VPWR _11976_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14663_ _14663_/A VGND VGND VPWR VPWR _15349_/A sky130_fd_sc_hd__buf_1
X_11875_ _11845_/X _11874_/Y _11845_/X _11874_/Y VGND VGND VPWR VPWR _11907_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16402_ _16402_/A _16402_/B VGND VGND VPWR VPWR _16402_/X sky130_fd_sc_hd__or2_1
X_13614_ _10428_/X _13613_/X _10428_/X _13613_/X VGND VGND VPWR VPWR _13615_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10826_ _10826_/A VGND VGND VPWR VPWR _10826_/Y sky130_fd_sc_hd__clkinvlp_2
X_14594_ _15042_/A _12078_/Y _12002_/Y _14526_/X VGND VGND VPWR VPWR _14594_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16333_ _16290_/Y _16331_/X _16332_/Y VGND VGND VPWR VPWR _16333_/X sky130_fd_sc_hd__o21a_1
X_10757_ _11966_/A _10772_/B VGND VGND VPWR VPWR _10899_/A sky130_fd_sc_hd__and2_1
X_13545_ _15040_/A _13512_/B _13512_/Y VGND VGND VPWR VPWR _13545_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16264_ _16264_/A _16264_/B VGND VGND VPWR VPWR _16264_/Y sky130_fd_sc_hd__nand2_1
X_13476_ _13448_/X _13475_/X _13448_/X _13475_/X VGND VGND VPWR VPWR _13477_/B sky130_fd_sc_hd__a2bb2oi_1
X_10688_ _11994_/A _10814_/B _10687_/Y VGND VGND VPWR VPWR _10689_/A sky130_fd_sc_hd__o21ai_2
XFILLER_9_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15215_ _15216_/A _15216_/B VGND VGND VPWR VPWR _15268_/A sky130_fd_sc_hd__and2_1
X_12427_ _11612_/A _11694_/B _12425_/Y _12426_/Y VGND VGND VPWR VPWR _12427_/X sky130_fd_sc_hd__o22a_2
X_16195_ _16106_/A _15807_/B _15807_/Y VGND VGND VPWR VPWR _16196_/A sky130_fd_sc_hd__o21ai_1
XFILLER_126_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12358_ _14063_/A _12299_/B _12299_/Y _12249_/X VGND VGND VPWR VPWR _12358_/X sky130_fd_sc_hd__a2bb2o_1
X_15146_ _15146_/A _15146_/B VGND VGND VPWR VPWR _15146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12289_ _12289_/A _12362_/B VGND VGND VPWR VPWR _12289_/Y sky130_fd_sc_hd__nand2_1
X_15077_ _15031_/X _15076_/X _15031_/X _15076_/X VGND VGND VPWR VPWR _15078_/B sky130_fd_sc_hd__a2bb2o_1
X_11309_ _11309_/A _11309_/B VGND VGND VPWR VPWR _11309_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14028_ _14028_/A VGND VGND VPWR VPWR _15461_/A sky130_fd_sc_hd__buf_1
XFILLER_122_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15979_ _15909_/Y _15978_/Y _15912_/Y VGND VGND VPWR VPWR _15979_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08520_ _09476_/B VGND VGND VPWR VPWR _08694_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08451_ _08710_/A VGND VGND VPWR VPWR _09331_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08382_ _08366_/A _08365_/Y _08366_/Y _08365_/A _08419_/A VGND VGND VPWR VPWR _08642_/A
+ sky130_fd_sc_hd__o221a_1
X_09003_ _11572_/A _09003_/B VGND VGND VPWR VPWR _12302_/A sky130_fd_sc_hd__or2_1
XFILLER_3_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09905_ _09857_/A _09857_/B _09904_/Y VGND VGND VPWR VPWR _10656_/A sky130_fd_sc_hd__a21oi_1
XFILLER_86_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _09836_/A VGND VGND VPWR VPWR _09836_/Y sky130_fd_sc_hd__inv_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09767_ _09730_/A _09730_/B _09733_/A VGND VGND VPWR VPWR _10052_/A sky130_fd_sc_hd__a21bo_1
XFILLER_67_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08718_ _08718_/A _09462_/B VGND VGND VPWR VPWR _08718_/Y sky130_fd_sc_hd__nor2_1
X_09698_ _09698_/A _09698_/B VGND VGND VPWR VPWR _09730_/A sky130_fd_sc_hd__or2_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08649_ input2/X input18/X _08392_/Y _08481_/Y _08392_/A VGND VGND VPWR VPWR _08650_/B
+ sky130_fd_sc_hd__o32a_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer50 _08667_/A VGND VGND VPWR VPWR _09679_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _12789_/A _11661_/B VGND VGND VPWR VPWR _11662_/A sky130_fd_sc_hd__and2_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11591_ _09429_/A _11591_/A2 _09750_/Y VGND VGND VPWR VPWR _11591_/Y sky130_fd_sc_hd__a21oi_1
X_10611_ _09954_/Y _10610_/A _09954_/A _10610_/Y _09797_/A VGND VGND VPWR VPWR _11888_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13330_ _13287_/A _13329_/Y _13287_/A _13329_/Y VGND VGND VPWR VPWR _13331_/B sky130_fd_sc_hd__a2bb2o_1
X_10542_ _09274_/A _09274_/B _09274_/X VGND VGND VPWR VPWR _10543_/B sky130_fd_sc_hd__a21boi_1
XFILLER_10_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13261_ _13925_/A VGND VGND VPWR VPWR _14724_/A sky130_fd_sc_hd__inv_2
XFILLER_41_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12212_ _12212_/A _12151_/X VGND VGND VPWR VPWR _12212_/X sky130_fd_sc_hd__or2b_1
X_15000_ _11752_/X _14999_/X _11754_/B VGND VGND VPWR VPWR _15000_/X sky130_fd_sc_hd__o21a_1
X_10473_ _11855_/A VGND VGND VPWR VPWR _12697_/A sky130_fd_sc_hd__buf_1
XFILLER_6_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13192_ _13192_/A _13192_/B VGND VGND VPWR VPWR _13192_/Y sky130_fd_sc_hd__nand2_1
X_12143_ _13921_/A _12143_/B VGND VGND VPWR VPWR _12143_/X sky130_fd_sc_hd__or2_1
X_12074_ _12073_/Y _11984_/X _12007_/Y VGND VGND VPWR VPWR _12074_/X sky130_fd_sc_hd__o21a_1
XFILLER_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15902_ _15902_/A _15902_/B VGND VGND VPWR VPWR _15902_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11025_ _12849_/A VGND VGND VPWR VPWR _15069_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15833_ _16192_/A VGND VGND VPWR VPWR _16160_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15764_ _14908_/A _14908_/B _14908_/Y VGND VGND VPWR VPWR _15764_/X sky130_fd_sc_hd__o21a_1
X_14715_ _14715_/A _14645_/X VGND VGND VPWR VPWR _14715_/X sky130_fd_sc_hd__or2b_1
X_12976_ _13698_/A VGND VGND VPWR VPWR _14411_/A sky130_fd_sc_hd__inv_2
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15695_ _15689_/Y _15693_/Y _15694_/Y VGND VGND VPWR VPWR _15695_/X sky130_fd_sc_hd__o21a_1
XFILLER_73_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11927_ _11928_/A _11928_/B VGND VGND VPWR VPWR _11927_/X sky130_fd_sc_hd__and2_1
X_14646_ _14715_/A _14644_/Y _14645_/X VGND VGND VPWR VPWR _14646_/Y sky130_fd_sc_hd__o21ai_1
X_11858_ _10458_/A _11810_/A _10556_/B _11857_/Y VGND VGND VPWR VPWR _11859_/A sky130_fd_sc_hd__o22a_1
XFILLER_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14577_ _14577_/A _14577_/B VGND VGND VPWR VPWR _14577_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11789_ _11722_/B _11788_/X _11722_/B _11788_/X VGND VGND VPWR VPWR _11790_/B sky130_fd_sc_hd__a2bb2o_1
X_10809_ _11990_/A VGND VGND VPWR VPWR _13509_/A sky130_fd_sc_hd__buf_1
XFILLER_13_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16316_ _16316_/A _16316_/B VGND VGND VPWR VPWR _16316_/Y sky130_fd_sc_hd__nand2_1
X_13528_ _10336_/Y _13480_/A _10336_/Y _13480_/A VGND VGND VPWR VPWR _13529_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16247_ _16241_/A _16246_/A _16241_/Y _16246_/Y _16238_/A VGND VGND VPWR VPWR _16248_/B
+ sky130_fd_sc_hd__a221o_1
X_13459_ _15171_/A VGND VGND VPWR VPWR _15425_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16178_ _16264_/A _16330_/A VGND VGND VPWR VPWR _16178_/Y sky130_fd_sc_hd__nor2_1
X_15129_ _15072_/A _15072_/B _15072_/Y VGND VGND VPWR VPWR _15129_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09621_ _09972_/A VGND VGND VPWR VPWR _09960_/A sky130_fd_sc_hd__buf_1
X_09552_ _09607_/A _09550_/X _09607_/B VGND VGND VPWR VPWR _09552_/X sky130_fd_sc_hd__o21ba_1
XFILLER_83_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08503_ _08701_/A _08503_/B VGND VGND VPWR VPWR _09448_/B sky130_fd_sc_hd__or2_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09483_ _08765_/A _09475_/X _08765_/A _09475_/X VGND VGND VPWR VPWR _09484_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_51_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08434_ _08434_/A VGND VGND VPWR VPWR _08434_/Y sky130_fd_sc_hd__inv_2
X_08365_ _08365_/A VGND VGND VPWR VPWR _08365_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08296_ _08296_/A VGND VGND VPWR VPWR _08296_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09819_ _09819_/A _09819_/B VGND VGND VPWR VPWR _09820_/B sky130_fd_sc_hd__or2_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _12830_/A _12830_/B VGND VGND VPWR VPWR _12830_/Y sky130_fd_sc_hd__nor2_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12761_ _12764_/A _12764_/B VGND VGND VPWR VPWR _12761_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _14794_/A _15455_/B _15455_/X _15479_/Y VGND VGND VPWR VPWR _15480_/X sky130_fd_sc_hd__o22a_1
X_11712_ _12065_/A VGND VGND VPWR VPWR _13198_/A sky130_fd_sc_hd__buf_1
X_14500_ _14500_/A VGND VGND VPWR VPWR _15211_/A sky130_fd_sc_hd__buf_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _10689_/A _12667_/A _10689_/Y _12667_/Y VGND VGND VPWR VPWR _12693_/B sky130_fd_sc_hd__o22a_1
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _13274_/A _14428_/B _14428_/Y _14430_/X VGND VGND VPWR VPWR _14431_/X sky130_fd_sc_hd__o2bb2a_1
X_11643_ _11640_/X _11642_/X _11640_/X _11642_/X VGND VGND VPWR VPWR _11644_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 wbs_dat_i[4] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__buf_4
XFILLER_128_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14362_ _11709_/A _14247_/A _14248_/B VGND VGND VPWR VPWR _15777_/A sky130_fd_sc_hd__o21ai_2
X_16101_ _16101_/A _16104_/B VGND VGND VPWR VPWR _16101_/Y sky130_fd_sc_hd__nor2_1
X_11574_ _12496_/A VGND VGND VPWR VPWR _15554_/A sky130_fd_sc_hd__buf_1
Xinput17 wbs_adr_i[9] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14293_ _14308_/A _14293_/B VGND VGND VPWR VPWR _15972_/A sky130_fd_sc_hd__or2_1
X_13313_ _13313_/A _13313_/B VGND VGND VPWR VPWR _13313_/X sky130_fd_sc_hd__and2_1
X_10525_ _11838_/A _10525_/B VGND VGND VPWR VPWR _10525_/Y sky130_fd_sc_hd__nand2_1
X_16032_ _16032_/A _16032_/B VGND VGND VPWR VPWR _16032_/Y sky130_fd_sc_hd__nand2_1
X_13244_ _13193_/X _13243_/Y _13193_/X _13243_/Y VGND VGND VPWR VPWR _13288_/B sky130_fd_sc_hd__a2bb2o_1
X_10456_ _09122_/A _10455_/X _09122_/A _10455_/X VGND VGND VPWR VPWR _11214_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13175_ _13184_/A VGND VGND VPWR VPWR _15331_/A sky130_fd_sc_hd__buf_1
XFILLER_6_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12126_ _12054_/X _12125_/Y _12054_/X _12125_/Y VGND VGND VPWR VPWR _12143_/B sky130_fd_sc_hd__a2bb2o_1
X_10387_ _10450_/A _11806_/A VGND VGND VPWR VPWR _10387_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12057_ _12057_/A _12057_/B VGND VGND VPWR VPWR _12057_/Y sky130_fd_sc_hd__nand2_1
X_11008_ _13897_/A _11094_/B VGND VGND VPWR VPWR _11186_/A sky130_fd_sc_hd__and2_1
X_15816_ _15731_/Y _15814_/X _15815_/Y VGND VGND VPWR VPWR _15816_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15747_ _15677_/A _15677_/B _15677_/Y VGND VGND VPWR VPWR _15747_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12959_ _14836_/A _13035_/B VGND VGND VPWR VPWR _13040_/A sky130_fd_sc_hd__and2_1
XFILLER_33_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15678_ _15614_/Y _15676_/X _15677_/Y VGND VGND VPWR VPWR _15678_/X sky130_fd_sc_hd__o21a_1
X_14629_ _15337_/A _14651_/B VGND VGND VPWR VPWR _14629_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08983_ _08880_/X _08981_/X _09001_/B VGND VGND VPWR VPWR _08983_/X sky130_fd_sc_hd__o21a_2
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09604_ _09494_/A _09494_/B _09494_/Y VGND VGND VPWR VPWR _09604_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09535_ _09551_/A _09551_/B VGND VGND VPWR VPWR _09607_/A sky130_fd_sc_hd__nor2_1
X_09466_ _10015_/A _08597_/A _09455_/Y _09465_/X VGND VGND VPWR VPWR _09466_/X sky130_fd_sc_hd__o22a_1
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08417_ _08351_/Y _08413_/Y _10016_/A VGND VGND VPWR VPWR _08417_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09397_ _12855_/A VGND VGND VPWR VPWR _15060_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08348_ _08348_/A VGND VGND VPWR VPWR _08348_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08279_ input9/X _08279_/B VGND VGND VPWR VPWR _08279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11290_ _12256_/A _11290_/B VGND VGND VPWR VPWR _11290_/Y sky130_fd_sc_hd__nor2_1
X_10310_ _10310_/A VGND VGND VPWR VPWR _10310_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10241_ _10241_/A _10241_/B VGND VGND VPWR VPWR _10241_/X sky130_fd_sc_hd__or2_1
X_10172_ _10124_/A _10124_/B _10125_/B VGND VGND VPWR VPWR _10173_/B sky130_fd_sc_hd__a21bo_1
XFILLER_121_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14980_ _15425_/A _14980_/B VGND VGND VPWR VPWR _14980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13931_ _15392_/A _13939_/B VGND VGND VPWR VPWR _14040_/A sky130_fd_sc_hd__and2_1
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13862_ _13776_/X _13791_/X _13793_/B VGND VGND VPWR VPWR _13862_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15601_ _15601_/A VGND VGND VPWR VPWR _15601_/Y sky130_fd_sc_hd__inv_2
X_13793_ _13791_/X _13793_/B VGND VGND VPWR VPWR _13793_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_62_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12813_ _12771_/X _12812_/Y _12771_/X _12812_/Y VGND VGND VPWR VPWR _12847_/B sky130_fd_sc_hd__a2bb2o_1
X_15532_ _14798_/A _15458_/B _15458_/Y VGND VGND VPWR VPWR _15532_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12714_/X _12743_/X _12714_/X _12743_/X VGND VGND VPWR VPWR _12774_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15463_ _15401_/X _15462_/X _15401_/X _15462_/X VGND VGND VPWR VPWR _15464_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12675_/A VGND VGND VPWR VPWR _12675_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15394_ _12045_/A _15393_/Y _12045_/A _15393_/Y VGND VGND VPWR VPWR _15396_/B sky130_fd_sc_hd__a2bb2o_1
X_14414_ _11788_/A _14413_/X _11787_/X VGND VGND VPWR VPWR _14415_/A sky130_fd_sc_hd__o21ai_2
X_11626_ _11626_/A VGND VGND VPWR VPWR _11627_/B sky130_fd_sc_hd__inv_2
X_14345_ _13419_/Y _14344_/X _13419_/Y _14344_/X VGND VGND VPWR VPWR _14346_/B sky130_fd_sc_hd__a2bb2oi_1
X_11557_ _14832_/A _11557_/B VGND VGND VPWR VPWR _11557_/X sky130_fd_sc_hd__or2_1
XFILLER_128_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10508_ _09836_/Y _10507_/Y _09836_/A _10507_/A _09941_/A VGND VGND VPWR VPWR _13608_/A
+ sky130_fd_sc_hd__o221a_2
X_16015_ _15953_/X _16014_/Y _15953_/X _16014_/Y VGND VGND VPWR VPWR _16036_/B sky130_fd_sc_hd__a2bb2o_1
X_14276_ _14276_/A VGND VGND VPWR VPWR _14276_/Y sky130_fd_sc_hd__inv_2
X_11488_ _12289_/A _11346_/B _11346_/Y _11285_/X VGND VGND VPWR VPWR _11488_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13227_ _14596_/A VGND VGND VPWR VPWR _14738_/A sky130_fd_sc_hd__buf_1
X_10439_ _10437_/A _10438_/A _10437_/Y _10438_/Y _09392_/A VGND VGND VPWR VPWR _10440_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13158_ _13114_/X _13157_/Y _13114_/X _13157_/Y VGND VGND VPWR VPWR _13196_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12109_ _13897_/A _12155_/B VGND VGND VPWR VPWR _12206_/A sky130_fd_sc_hd__and2_1
XFILLER_85_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13089_ _13758_/A VGND VGND VPWR VPWR _15264_/A sky130_fd_sc_hd__buf_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09320_ _09470_/B _09859_/A _09353_/A VGND VGND VPWR VPWR _09320_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09251_ _09251_/A _09251_/B VGND VGND VPWR VPWR _10065_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09182_ _09430_/A _09185_/B VGND VGND VPWR VPWR _09182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08966_ _09547_/A _08622_/A _08624_/A VGND VGND VPWR VPWR _08966_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08897_ _09553_/A _08584_/A _08586_/A VGND VGND VPWR VPWR _08897_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09518_ _09518_/A _09518_/B VGND VGND VPWR VPWR _09518_/X sky130_fd_sc_hd__and2_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10790_ _12070_/A VGND VGND VPWR VPWR _13700_/A sky130_fd_sc_hd__buf_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09449_ _09482_/A _09525_/A VGND VGND VPWR VPWR _09449_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12460_ _13882_/A _12460_/B VGND VGND VPWR VPWR _12460_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11411_ _11413_/A _11411_/B VGND VGND VPWR VPWR _12322_/A sky130_fd_sc_hd__or2_1
X_12391_ _13974_/A _12451_/B _12390_/Y VGND VGND VPWR VPWR _12391_/Y sky130_fd_sc_hd__o21ai_1
X_14130_ _14131_/A _14132_/A VGND VGND VPWR VPWR _14130_/Y sky130_fd_sc_hd__nor2_1
X_11342_ _11298_/X _11341_/Y _11298_/X _11341_/Y VGND VGND VPWR VPWR _11493_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14061_ _14061_/A _14061_/B VGND VGND VPWR VPWR _14128_/B sky130_fd_sc_hd__or2_1
X_11273_ _11506_/A VGND VGND VPWR VPWR _13785_/A sky130_fd_sc_hd__buf_1
XFILLER_79_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13012_ _13676_/A _13012_/B VGND VGND VPWR VPWR _13012_/Y sky130_fd_sc_hd__nand2_1
X_10224_ _10224_/A _10224_/B VGND VGND VPWR VPWR _10309_/A sky130_fd_sc_hd__and2_1
XFILLER_4_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10155_ _10155_/A _10155_/B VGND VGND VPWR VPWR _10155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14963_ _14933_/Y _14962_/Y _14933_/Y _14962_/Y VGND VGND VPWR VPWR _14982_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10086_ _10040_/X _10084_/X _11318_/B VGND VGND VPWR VPWR _10086_/X sky130_fd_sc_hd__o21a_1
X_14894_ _14818_/X _14893_/X _14818_/X _14893_/X VGND VGND VPWR VPWR _14910_/B sky130_fd_sc_hd__a2bb2o_1
X_13914_ _14622_/A _13847_/B _13847_/Y VGND VGND VPWR VPWR _13914_/Y sky130_fd_sc_hd__o21ai_1
X_13845_ _14626_/A _13845_/B VGND VGND VPWR VPWR _13845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13776_ _13703_/X _13718_/X _13720_/B VGND VGND VPWR VPWR _13776_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10988_ _11138_/A _12689_/A _10987_/Y VGND VGND VPWR VPWR _10988_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15515_ _15512_/A _15512_/B _15512_/X _15651_/A VGND VGND VPWR VPWR _15519_/B sky130_fd_sc_hd__o22a_1
X_12727_ _12786_/A _12786_/B VGND VGND VPWR VPWR _12727_/Y sky130_fd_sc_hd__nor2_1
X_15446_ _15446_/A _15446_/B VGND VGND VPWR VPWR _15446_/X sky130_fd_sc_hd__and2_1
X_12658_ _10201_/Y _12657_/Y _10213_/Y VGND VGND VPWR VPWR _12658_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_128_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11609_ _10194_/A _11609_/A2 _10194_/Y VGND VGND VPWR VPWR _11610_/A sky130_fd_sc_hd__o21ai_1
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12589_ _12586_/Y _12588_/Y _12586_/A _12588_/A _11708_/A VGND VGND VPWR VPWR _12620_/A
+ sky130_fd_sc_hd__o221a_1
X_15377_ _15408_/A _15408_/B VGND VGND VPWR VPWR _15453_/A sky130_fd_sc_hd__and2_1
X_14328_ _14334_/A _14328_/B VGND VGND VPWR VPWR _15958_/A sky130_fd_sc_hd__or2_1
X_14259_ _15872_/A _14259_/B VGND VGND VPWR VPWR _14259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _09251_/A VGND VGND VPWR VPWR _09498_/A sky130_fd_sc_hd__buf_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _09338_/B VGND VGND VPWR VPWR _10134_/A sky130_fd_sc_hd__buf_1
XFILLER_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08682_ _09538_/A _08635_/A _08637_/Y _08681_/Y VGND VGND VPWR VPWR _08682_/X sky130_fd_sc_hd__o22a_1
XFILLER_66_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09303_ _09303_/A _10235_/A VGND VGND VPWR VPWR _09303_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09234_ _09234_/A _09681_/A VGND VGND VPWR VPWR _09629_/A sky130_fd_sc_hd__or2_1
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09165_ _10010_/B _09165_/B VGND VGND VPWR VPWR _09166_/B sky130_fd_sc_hd__or2_1
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09096_ _09716_/A VGND VGND VPWR VPWR _09717_/A sky130_fd_sc_hd__buf_1
XFILLER_102_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09998_ _09964_/X _11513_/A _11512_/B VGND VGND VPWR VPWR _09999_/B sky130_fd_sc_hd__o21ai_1
XFILLER_130_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08949_ _09459_/B VGND VGND VPWR VPWR _09539_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11960_ _11966_/A _11966_/B VGND VGND VPWR VPWR _12040_/A sky130_fd_sc_hd__and2_1
XFILLER_57_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10911_ _13832_/A _10910_/B _11067_/A _10910_/Y VGND VGND VPWR VPWR _10911_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11891_ _10626_/A _11890_/X _10626_/A _11890_/X VGND VGND VPWR VPWR _11893_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10842_ _12070_/A _10938_/B VGND VGND VPWR VPWR _10842_/Y sky130_fd_sc_hd__nand2_1
X_13630_ _13595_/Y _13627_/Y _13629_/Y VGND VGND VPWR VPWR _13631_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10773_ _10899_/A _10770_/X _10772_/X VGND VGND VPWR VPWR _10773_/X sky130_fd_sc_hd__o21a_1
X_13561_ _15032_/A _13524_/B _13524_/Y VGND VGND VPWR VPWR _13561_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16280_ _16271_/X _16279_/Y _16271_/X _16279_/Y VGND VGND VPWR VPWR _16338_/B sky130_fd_sc_hd__o2bb2a_1
X_12512_ _12511_/A _12511_/B _12511_/Y _12503_/X VGND VGND VPWR VPWR _12638_/B sky130_fd_sc_hd__o211a_1
X_15300_ _14664_/A _15243_/B _15243_/Y VGND VGND VPWR VPWR _15300_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15231_ _15285_/A _15285_/B VGND VGND VPWR VPWR _15287_/A sky130_fd_sc_hd__nor2_1
X_13492_ _11621_/Y _12382_/A _11538_/Y _13491_/X VGND VGND VPWR VPWR _13492_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12443_ _13871_/A _12442_/B _12442_/X _12370_/X VGND VGND VPWR VPWR _12443_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12374_ _13495_/A VGND VGND VPWR VPWR _12437_/A sky130_fd_sc_hd__clkinvlp_2
X_15162_ _12422_/A _15161_/Y _12422_/A _15161_/Y VGND VGND VPWR VPWR _15163_/B sky130_fd_sc_hd__a2bb2o_1
X_14113_ _14113_/A VGND VGND VPWR VPWR _14880_/A sky130_fd_sc_hd__inv_2
XFILLER_99_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15093_ _15072_/A _15072_/B _15072_/Y _15092_/X VGND VGND VPWR VPWR _15093_/X sky130_fd_sc_hd__a2bb2o_1
X_11325_ _11325_/A1 _11323_/Y _11324_/Y _11323_/A _11529_/A VGND VGND VPWR VPWR _11521_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11256_ _14035_/A _11231_/B _11231_/Y _11255_/X VGND VGND VPWR VPWR _11256_/X sky130_fd_sc_hd__a2bb2o_1
X_14044_ _14429_/A _13937_/B _14429_/A _13937_/B VGND VGND VPWR VPWR _14044_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11187_ _11093_/X _11186_/X _11093_/X _11186_/X VGND VGND VPWR VPWR _11188_/B sky130_fd_sc_hd__a2bb2o_1
X_10207_ _10346_/B VGND VGND VPWR VPWR _10462_/A sky130_fd_sc_hd__clkbuf_2
X_15995_ _16055_/A _16055_/B VGND VGND VPWR VPWR _15995_/X sky130_fd_sc_hd__and2_1
XFILLER_95_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10138_ _10133_/A _10133_/B _10134_/B VGND VGND VPWR VPWR _10139_/B sky130_fd_sc_hd__a21bo_1
X_14946_ _14943_/Y _14945_/X _14943_/Y _14945_/X VGND VGND VPWR VPWR _14948_/B sky130_fd_sc_hd__a2bb2o_1
X_10069_ _10069_/A _10069_/B VGND VGND VPWR VPWR _10069_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14877_ _14786_/A _14786_/B _14786_/A _14786_/B VGND VGND VPWR VPWR _14877_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13828_ _13828_/A VGND VGND VPWR VPWR _14645_/A sky130_fd_sc_hd__inv_2
X_13759_ _13825_/A _13757_/X _13758_/X VGND VGND VPWR VPWR _13759_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15429_ _15424_/Y _15428_/X _15424_/Y _15428_/X VGND VGND VPWR VPWR _15429_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09921_ _09918_/X _09921_/B VGND VGND VPWR VPWR _09923_/B sky130_fd_sc_hd__nand2b_1
XFILLER_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09852_ _09853_/A _09853_/B VGND VGND VPWR VPWR _09855_/A sky130_fd_sc_hd__nor2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _10014_/A _10128_/A VGND VGND VPWR VPWR _08803_/Y sky130_fd_sc_hd__nor2_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _10083_/A _09781_/Y _09782_/Y VGND VGND VPWR VPWR _09785_/B sky130_fd_sc_hd__o21ai_1
XFILLER_100_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08734_ _10012_/A _09531_/A VGND VGND VPWR VPWR _08734_/X sky130_fd_sc_hd__or2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08665_ _08665_/A VGND VGND VPWR VPWR _08671_/A sky130_fd_sc_hd__inv_2
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08596_ _08596_/A VGND VGND VPWR VPWR _10114_/B sky130_fd_sc_hd__inv_2
XFILLER_41_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09217_ _09217_/A _09217_/B VGND VGND VPWR VPWR _09803_/A sky130_fd_sc_hd__or2_2
X_09148_ _08762_/A _09147_/X _08532_/B VGND VGND VPWR VPWR _09148_/X sky130_fd_sc_hd__o21ba_1
XFILLER_108_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09079_ _10011_/B _09078_/B _09165_/B VGND VGND VPWR VPWR _09760_/A sky130_fd_sc_hd__a21bo_1
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ _12103_/A _11000_/B _11000_/Y _10932_/X VGND VGND VPWR VPWR _11110_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12090_ _12090_/A _12089_/X VGND VGND VPWR VPWR _12090_/X sky130_fd_sc_hd__or2b_1
X_11041_ _13917_/A _11084_/B VGND VGND VPWR VPWR _11223_/A sky130_fd_sc_hd__and2_1
XFILLER_1_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14800_ _14800_/A _14728_/X VGND VGND VPWR VPWR _14800_/X sky130_fd_sc_hd__or2b_1
XFILLER_76_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15780_ _15785_/A _15785_/B VGND VGND VPWR VPWR _16245_/A sky130_fd_sc_hd__and2_1
XFILLER_85_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12992_ _12992_/A VGND VGND VPWR VPWR _13672_/A sky130_fd_sc_hd__inv_2
X_14731_ _14796_/A _14729_/X _14730_/X VGND VGND VPWR VPWR _14731_/X sky130_fd_sc_hd__o21a_1
X_11943_ _13696_/A _11910_/B _11910_/Y VGND VGND VPWR VPWR _11943_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14662_ _14609_/Y _14660_/X _14661_/Y VGND VGND VPWR VPWR _14662_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11874_ _11846_/A _11846_/B _11846_/Y VGND VGND VPWR VPWR _11874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16401_ _16394_/Y _16398_/Y _16399_/Y _16400_/Y VGND VGND VPWR VPWR _16401_/X sky130_fd_sc_hd__o211a_1
X_13613_ _12915_/A _14429_/B _12915_/A _14429_/B VGND VGND VPWR VPWR _13613_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10825_ _12084_/A _10966_/B _10824_/Y VGND VGND VPWR VPWR _10826_/A sky130_fd_sc_hd__o21ai_2
X_16332_ _16332_/A _16332_/B VGND VGND VPWR VPWR _16332_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14593_ _14528_/A _14528_/B _14525_/X _14528_/Y VGND VGND VPWR VPWR _14593_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13544_ _13544_/A VGND VGND VPWR VPWR _15420_/A sky130_fd_sc_hd__buf_1
X_10756_ _10630_/X _10755_/Y _10630_/X _10755_/Y VGND VGND VPWR VPWR _10772_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16263_ _16186_/Y _16261_/X _16262_/Y VGND VGND VPWR VPWR _16263_/X sky130_fd_sc_hd__o21a_1
X_13475_ _13449_/A _13449_/B _13449_/Y VGND VGND VPWR VPWR _13475_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10687_ _11994_/A _10814_/B VGND VGND VPWR VPWR _10687_/Y sky130_fd_sc_hd__nand2_1
X_16194_ _16260_/A _16326_/A VGND VGND VPWR VPWR _16194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15214_ _10522_/Y _15213_/Y _10522_/Y _15213_/Y VGND VGND VPWR VPWR _15216_/B sky130_fd_sc_hd__o2bb2a_1
X_12426_ _12426_/A _12426_/B VGND VGND VPWR VPWR _12426_/Y sky130_fd_sc_hd__nor2_1
X_15145_ _12836_/X _15144_/X _12836_/X _15144_/X VGND VGND VPWR VPWR _15146_/B sky130_fd_sc_hd__a2bb2o_1
X_12357_ _12302_/A _12302_/B _12302_/Y _12511_/A VGND VGND VPWR VPWR _12412_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12288_ _12365_/A _12287_/Y _12365_/A _12287_/Y VGND VGND VPWR VPWR _12362_/B sky130_fd_sc_hd__a2bb2o_1
X_15076_ _15076_/A _15032_/X VGND VGND VPWR VPWR _15076_/X sky130_fd_sc_hd__or2b_1
X_11308_ _09965_/X _11308_/B VGND VGND VPWR VPWR _11309_/B sky130_fd_sc_hd__and2b_1
X_11239_ _11239_/A _11251_/B VGND VGND VPWR VPWR _14042_/A sky130_fd_sc_hd__or2_1
X_14027_ _14027_/A _14027_/B VGND VGND VPWR VPWR _14027_/X sky130_fd_sc_hd__and2_1
XFILLER_96_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15978_ _15978_/A _15978_/B VGND VGND VPWR VPWR _15978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14929_ _14863_/Y _14927_/X _14928_/Y VGND VGND VPWR VPWR _14929_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08450_ _10010_/A VGND VGND VPWR VPWR _08710_/A sky130_fd_sc_hd__inv_2
XFILLER_51_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08381_ _08401_/A VGND VGND VPWR VPWR _08419_/A sky130_fd_sc_hd__buf_6
XFILLER_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09002_ _08981_/X _09001_/X _08981_/X _09001_/X VGND VGND VPWR VPWR _09003_/B sky130_fd_sc_hd__a2bb2oi_4
XFILLER_117_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09904_ _09904_/A VGND VGND VPWR VPWR _09904_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09835_ _09799_/A _09799_/B _09834_/Y VGND VGND VPWR VPWR _09836_/A sky130_fd_sc_hd__a21oi_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09766_ _09766_/A VGND VGND VPWR VPWR _09776_/A sky130_fd_sc_hd__inv_2
XFILLER_66_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08717_ _08717_/A _08717_/B VGND VGND VPWR VPWR _08717_/X sky130_fd_sc_hd__or2_1
X_09697_ _08592_/A _09728_/B _08592_/A _09728_/B VGND VGND VPWR VPWR _09698_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer40 _08368_/X VGND VGND VPWR VPWR _08415_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer51 _08667_/A VGND VGND VPWR VPWR _10105_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_08648_ _09230_/A _10110_/B VGND VGND VPWR VPWR _08648_/X sky130_fd_sc_hd__or2_1
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08579_ _09209_/B VGND VGND VPWR VPWR _08579_/Y sky130_fd_sc_hd__inv_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11590_ _11590_/A _11590_/B VGND VGND VPWR VPWR _12445_/A sky130_fd_sc_hd__or2_2
X_10610_ _10610_/A VGND VGND VPWR VPWR _10610_/Y sky130_fd_sc_hd__inv_2
X_10541_ _13555_/A _10540_/B _10540_/X _10435_/X VGND VGND VPWR VPWR _10541_/X sky130_fd_sc_hd__o22a_1
XFILLER_127_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13260_ _14726_/A _13279_/B VGND VGND VPWR VPWR _13260_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12211_ _14017_/A _12211_/B VGND VGND VPWR VPWR _12211_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10472_ _10468_/Y _10470_/A _10468_/A _10470_/Y _10984_/A VGND VGND VPWR VPWR _11855_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_6_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13191_ _13168_/Y _13189_/X _13190_/Y VGND VGND VPWR VPWR _13191_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12142_ _12227_/A _12140_/X _12141_/X VGND VGND VPWR VPWR _12142_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12073_ _13640_/A _12073_/B VGND VGND VPWR VPWR _12073_/Y sky130_fd_sc_hd__nor2_1
X_15901_ _15862_/Y _15899_/X _15900_/Y VGND VGND VPWR VPWR _15901_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11024_ _13551_/A VGND VGND VPWR VPWR _12849_/A sky130_fd_sc_hd__buf_1
XFILLER_1_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15832_ _15832_/A VGND VGND VPWR VPWR _16192_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15763_ _16096_/A VGND VGND VPWR VPWR _16099_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12975_ _14523_/A _13027_/B VGND VGND VPWR VPWR _13060_/A sky130_fd_sc_hd__and2_1
X_14714_ _15392_/A VGND VGND VPWR VPWR _15398_/A sky130_fd_sc_hd__buf_1
XFILLER_80_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11926_ _10689_/A _11925_/A _10689_/Y _11994_/B VGND VGND VPWR VPWR _11928_/B sky130_fd_sc_hd__o22a_1
XFILLER_18_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15694_ _15694_/A _15694_/B VGND VGND VPWR VPWR _15694_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14645_ _14645_/A _14645_/B VGND VGND VPWR VPWR _14645_/X sky130_fd_sc_hd__or2_1
XFILLER_60_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11857_ _11857_/A _11857_/B VGND VGND VPWR VPWR _11857_/Y sky130_fd_sc_hd__nor2_1
X_14576_ _14562_/Y _14574_/X _14575_/Y VGND VGND VPWR VPWR _14576_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11788_ _11788_/A _11787_/X VGND VGND VPWR VPWR _11788_/X sky130_fd_sc_hd__or2b_1
XFILLER_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10808_ _10079_/A _10807_/Y _09968_/Y _10807_/A _10959_/A VGND VGND VPWR VPWR _11990_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16315_ _16316_/A _16316_/B VGND VGND VPWR VPWR _16315_/Y sky130_fd_sc_hd__nor2_1
X_10739_ _12992_/A _10639_/B _10639_/Y VGND VGND VPWR VPWR _10739_/Y sky130_fd_sc_hd__o21ai_1
X_13527_ _13527_/A _13527_/B VGND VGND VPWR VPWR _13527_/Y sky130_fd_sc_hd__nand2_1
X_16246_ _16246_/A VGND VGND VPWR VPWR _16246_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_9_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13458_ _13457_/Y _12787_/X _12723_/Y VGND VGND VPWR VPWR _13458_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16177_ _16264_/B VGND VGND VPWR VPWR _16330_/A sky130_fd_sc_hd__buf_6
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13389_ _14119_/A _13439_/B VGND VGND VPWR VPWR _13389_/Y sky130_fd_sc_hd__nor2_1
X_12409_ _12358_/X _12408_/Y _12358_/X _12408_/Y VGND VGND VPWR VPWR _12410_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15128_ _15128_/A _15128_/B VGND VGND VPWR VPWR _15128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15059_ _15043_/X _15058_/X _15043_/X _15058_/X VGND VGND VPWR VPWR _15060_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09620_ _09507_/X _09619_/X _09507_/X _09619_/X VGND VGND VPWR VPWR _09972_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09551_ _09551_/A _09551_/B VGND VGND VPWR VPWR _09607_/B sky130_fd_sc_hd__and2_1
X_08502_ _08308_/Y _08501_/A _08308_/A _08501_/Y VGND VGND VPWR VPWR _08503_/B sky130_fd_sc_hd__o22a_1
XFILLER_102_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09482_ _09482_/A _09482_/B VGND VGND VPWR VPWR _09482_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08433_ _09209_/B _08428_/X _09323_/A VGND VGND VPWR VPWR _08433_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08364_ _08364_/A _08364_/B VGND VGND VPWR VPWR _08365_/A sky130_fd_sc_hd__or2_1
XFILLER_11_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08295_ input22/X _08306_/B _08307_/A _08309_/A VGND VGND VPWR VPWR _08296_/A sky130_fd_sc_hd__o22a_1
XFILLER_117_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09818_ _09818_/A _09818_/B VGND VGND VPWR VPWR _09819_/B sky130_fd_sc_hd__or2_1
XFILLER_101_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09749_ _10034_/A VGND VGND VPWR VPWR _09749_/X sky130_fd_sc_hd__buf_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12760_ _12709_/X _12759_/X _12709_/X _12759_/X VGND VGND VPWR VPWR _12764_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11569_/A _11569_/B _11569_/Y _11710_/X VGND VGND VPWR VPWR _12640_/A sky130_fd_sc_hd__o211a_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12691_/A _12691_/B VGND VGND VPWR VPWR _12691_/Y sky130_fd_sc_hd__nor2_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _15396_/A _14429_/B _10428_/X _14429_/X VGND VGND VPWR VPWR _14430_/X sky130_fd_sc_hd__o22a_1
XFILLER_70_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11642_ _11641_/Y _11501_/X _11546_/Y VGND VGND VPWR VPWR _11642_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14361_ _14367_/A _14361_/B VGND VGND VPWR VPWR _14363_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16100_ _16096_/Y _16098_/X _16099_/Y VGND VGND VPWR VPWR _16104_/B sky130_fd_sc_hd__o21ai_1
X_11573_ _14148_/A VGND VGND VPWR VPWR _12496_/A sky130_fd_sc_hd__clkinvlp_2
X_13312_ _13305_/A _13311_/Y _13305_/A _13311_/Y VGND VGND VPWR VPWR _13313_/B sky130_fd_sc_hd__a2bb2o_1
Xinput18 wbs_dat_i[0] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_2
Xinput29 wbs_dat_i[5] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_4
XFILLER_109_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14292_ _13446_/X _14291_/X _13446_/X _14291_/X VGND VGND VPWR VPWR _14293_/B sky130_fd_sc_hd__a2bb2oi_1
X_10524_ _13609_/A _10523_/B _10522_/Y _10523_/Y VGND VGND VPWR VPWR _10524_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16031_ _16025_/Y _16029_/X _16030_/Y VGND VGND VPWR VPWR _16031_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13243_ _13194_/A _13194_/B _13194_/Y VGND VGND VPWR VPWR _13243_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10455_ _09418_/A _09123_/B _09123_/Y VGND VGND VPWR VPWR _10455_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13174_ _13824_/A _13186_/B VGND VGND VPWR VPWR _13174_/Y sky130_fd_sc_hd__nor2_1
X_12125_ _13188_/A _12055_/B _12055_/Y VGND VGND VPWR VPWR _12125_/Y sky130_fd_sc_hd__o21ai_1
X_10386_ _11806_/A VGND VGND VPWR VPWR _12699_/A sky130_fd_sc_hd__buf_1
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12056_ _12036_/Y _12054_/X _12055_/Y VGND VGND VPWR VPWR _12056_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11007_ _10926_/X _11006_/X _10926_/X _11006_/X VGND VGND VPWR VPWR _11094_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15815_ _16114_/A _15815_/B VGND VGND VPWR VPWR _15815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15746_ _15752_/A _15746_/B VGND VGND VPWR VPWR _16108_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12958_ _12947_/X _12957_/Y _12947_/X _12957_/Y VGND VGND VPWR VPWR _13035_/B sky130_fd_sc_hd__a2bb2o_1
X_15677_ _15677_/A _15677_/B VGND VGND VPWR VPWR _15677_/Y sky130_fd_sc_hd__nand2_1
X_11909_ _11909_/A VGND VGND VPWR VPWR _11909_/Y sky130_fd_sc_hd__inv_2
X_12889_ _12936_/A VGND VGND VPWR VPWR _14468_/A sky130_fd_sc_hd__buf_1
X_14628_ _14578_/X _14627_/Y _14578_/X _14627_/Y VGND VGND VPWR VPWR _14651_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14559_ _15264_/A VGND VGND VPWR VPWR _14575_/A sky130_fd_sc_hd__buf_1
XFILLER_9_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16229_ _16227_/A _16228_/A _16227_/Y _16228_/Y _15832_/A VGND VGND VPWR VPWR _16251_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08982_ _08982_/A _08982_/B VGND VGND VPWR VPWR _09001_/B sky130_fd_sc_hd__or2_1
XFILLER_130_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09603_ _09984_/A _09656_/B VGND VGND VPWR VPWR _09603_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09534_ _09553_/A _09553_/B VGND VGND VPWR VPWR _09601_/A sky130_fd_sc_hd__nor2_1
X_09465_ _10016_/A _08610_/A _09456_/Y _09464_/X VGND VGND VPWR VPWR _09465_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08416_ _09221_/A VGND VGND VPWR VPWR _10016_/A sky130_fd_sc_hd__buf_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09396_ _13648_/A VGND VGND VPWR VPWR _12855_/A sky130_fd_sc_hd__buf_1
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08347_ _08347_/A _08347_/B VGND VGND VPWR VPWR _08348_/A sky130_fd_sc_hd__or2_1
X_08278_ _08278_/A VGND VGND VPWR VPWR _08279_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10240_ _10240_/A _10240_/B VGND VGND VPWR VPWR _10240_/X sky130_fd_sc_hd__or2_1
XFILLER_133_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10171_ _10111_/A _10111_/B _10112_/A VGND VGND VPWR VPWR _10173_/A sky130_fd_sc_hd__a21bo_1
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13930_ _13838_/X _13929_/Y _13838_/X _13929_/Y VGND VGND VPWR VPWR _13939_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15600_ _15600_/A _15542_/X VGND VGND VPWR VPWR _15601_/A sky130_fd_sc_hd__or2b_1
X_13861_ _13775_/X _13795_/X _13797_/B VGND VGND VPWR VPWR _13861_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13792_ _13792_/A _13792_/B VGND VGND VPWR VPWR _13793_/B sky130_fd_sc_hd__or2_1
X_12812_ _12772_/A _12772_/B _12772_/Y VGND VGND VPWR VPWR _12812_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15531_ _15534_/A _15534_/B VGND VGND VPWR VPWR _15531_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12695_/A _12695_/B _12695_/Y VGND VGND VPWR VPWR _12743_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15462_ _15462_/A _15402_/X VGND VGND VPWR VPWR _15462_/X sky130_fd_sc_hd__or2b_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _12833_/A _11720_/B _14412_/X VGND VGND VPWR VPWR _14413_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12674_ _11316_/Y _12673_/Y _11150_/Y VGND VGND VPWR VPWR _12675_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15393_ _15329_/A _15329_/B _15329_/Y VGND VGND VPWR VPWR _15393_/Y sky130_fd_sc_hd__a21oi_1
X_11625_ _11620_/Y _11624_/Y _11620_/Y _11624_/Y VGND VGND VPWR VPWR _11626_/A sky130_fd_sc_hd__a2bb2o_1
X_14344_ _14095_/A _13420_/B _13420_/Y VGND VGND VPWR VPWR _14344_/X sky130_fd_sc_hd__o21a_1
X_11556_ _12400_/A VGND VGND VPWR VPWR _14832_/A sky130_fd_sc_hd__buf_1
XFILLER_11_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14275_ _14185_/Y _14273_/Y _14274_/Y VGND VGND VPWR VPWR _14275_/Y sky130_fd_sc_hd__o21ai_1
X_10507_ _10507_/A VGND VGND VPWR VPWR _10507_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16014_ _15936_/X _16014_/B VGND VGND VPWR VPWR _16014_/Y sky130_fd_sc_hd__nand2b_1
X_13226_ _15060_/A VGND VGND VPWR VPWR _14596_/A sky130_fd_sc_hd__inv_2
X_11487_ _13206_/A VGND VGND VPWR VPWR _12400_/A sky130_fd_sc_hd__clkinvlp_2
X_10438_ _10438_/A VGND VGND VPWR VPWR _10438_/Y sky130_fd_sc_hd__inv_2
X_13157_ _15249_/A _13115_/B _13115_/Y VGND VGND VPWR VPWR _13157_/Y sky130_fd_sc_hd__o21ai_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _11762_/A _10369_/B VGND VGND VPWR VPWR _10369_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12108_ _12066_/X _12107_/Y _12066_/X _12107_/Y VGND VGND VPWR VPWR _12155_/B sky130_fd_sc_hd__a2bb2o_1
X_13088_ _13088_/A VGND VGND VPWR VPWR _13758_/A sky130_fd_sc_hd__inv_2
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12039_ _12039_/A _12053_/B VGND VGND VPWR VPWR _12039_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15729_ _15683_/A _15683_/B _15683_/Y VGND VGND VPWR VPWR _15729_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09250_ _09456_/A _09250_/B VGND VGND VPWR VPWR _10069_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09181_ _09177_/Y _09179_/Y _09180_/Y VGND VGND VPWR VPWR _09185_/B sky130_fd_sc_hd__o21ai_1
XFILLER_107_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08965_ _08968_/A _08968_/B VGND VGND VPWR VPWR _08965_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08896_ _08976_/A _08976_/B VGND VGND VPWR VPWR _08896_/X sky130_fd_sc_hd__and2_1
XFILLER_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09517_ _09482_/A _09482_/B _09482_/Y _09516_/X VGND VGND VPWR VPWR _09563_/A sky130_fd_sc_hd__o2bb2a_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _09448_/A _09448_/B VGND VGND VPWR VPWR _09448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09379_ _09379_/A VGND VGND VPWR VPWR _09432_/B sky130_fd_sc_hd__inv_2
X_12390_ _12390_/A _12451_/B VGND VGND VPWR VPWR _12390_/Y sky130_fd_sc_hd__nand2_1
X_11410_ _11407_/Y _11409_/Y _11407_/A _11409_/A _12606_/B VGND VGND VPWR VPWR _14083_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11341_ _13788_/A _11500_/B _11340_/Y VGND VGND VPWR VPWR _11341_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14060_ _14122_/A _14058_/X _14059_/X VGND VGND VPWR VPWR _14060_/X sky130_fd_sc_hd__o21a_1
X_11272_ _11271_/A _11271_/B _11271_/Y _09392_/X VGND VGND VPWR VPWR _11506_/A sky130_fd_sc_hd__o211a_1
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13011_ _14504_/A _13010_/B _13009_/Y _13010_/Y VGND VGND VPWR VPWR _13011_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10223_ _10175_/Y _10222_/A _10175_/A _10222_/Y _10462_/A VGND VGND VPWR VPWR _10224_/B
+ sky130_fd_sc_hd__a221o_1
X_10154_ _08793_/B _10129_/B _10130_/B VGND VGND VPWR VPWR _10155_/B sky130_fd_sc_hd__a21bo_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14962_ _14971_/A _14971_/B _14961_/Y VGND VGND VPWR VPWR _14962_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10085_ _10085_/A _10085_/B VGND VGND VPWR VPWR _11318_/B sky130_fd_sc_hd__or2_1
X_14893_ _14806_/A _14806_/B _14806_/A _14806_/B VGND VGND VPWR VPWR _14893_/X sky130_fd_sc_hd__a2bb2o_1
X_13913_ _13913_/A VGND VGND VPWR VPWR _15406_/A sky130_fd_sc_hd__buf_1
XFILLER_90_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13844_ _13823_/Y _13842_/X _13843_/Y VGND VGND VPWR VPWR _13844_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13775_ _13722_/X _13773_/X _13800_/B VGND VGND VPWR VPWR _13775_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10987_ _11138_/A _12174_/A VGND VGND VPWR VPWR _10987_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15514_ _15474_/X _15513_/Y _15474_/X _15513_/Y VGND VGND VPWR VPWR _15651_/A sky130_fd_sc_hd__a2bb2o_1
X_12726_ _12720_/X _12725_/X _12720_/X _12725_/X VGND VGND VPWR VPWR _12786_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15445_ _15413_/X _15444_/X _15413_/X _15444_/X VGND VGND VPWR VPWR _15446_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12657_ _10282_/Y _12657_/A2 _10349_/A VGND VGND VPWR VPWR _12657_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15376_ _15340_/X _15375_/X _15340_/X _15375_/X VGND VGND VPWR VPWR _15408_/B sky130_fd_sc_hd__a2bb2o_1
X_11608_ _12426_/A VGND VGND VPWR VPWR _11612_/A sky130_fd_sc_hd__inv_2
X_12588_ _12588_/A VGND VGND VPWR VPWR _12588_/Y sky130_fd_sc_hd__inv_2
X_14327_ _13434_/Y _14326_/X _13434_/Y _14326_/X VGND VGND VPWR VPWR _14328_/B sky130_fd_sc_hd__a2bb2oi_1
X_11539_ _11623_/A _12419_/A _11538_/Y VGND VGND VPWR VPWR _11539_/X sky130_fd_sc_hd__a21o_1
X_14258_ _14258_/A VGND VGND VPWR VPWR _14258_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14189_ _14189_/A _12632_/X VGND VGND VPWR VPWR _14189_/X sky130_fd_sc_hd__or2b_1
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13209_ _14934_/A _13451_/B VGND VGND VPWR VPWR _13209_/Y sky130_fd_sc_hd__nand2_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08749_/A _08748_/Y _08749_/Y _09340_/B VGND VGND VPWR VPWR _09338_/B sky130_fd_sc_hd__o22a_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08681_ _09230_/A _10110_/B _08648_/X _08680_/X VGND VGND VPWR VPWR _08681_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09302_ _09303_/A _10235_/A VGND VGND VPWR VPWR _09302_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09233_ _09400_/A VGND VGND VPWR VPWR _09681_/A sky130_fd_sc_hd__inv_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09164_ _08765_/Y _09158_/A _08765_/A _09158_/Y VGND VGND VPWR VPWR _10010_/B sky130_fd_sc_hd__o22a_1
XFILLER_119_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09095_ _10018_/B _09071_/B _09072_/B VGND VGND VPWR VPWR _09716_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09997_ _09997_/A _09997_/B VGND VGND VPWR VPWR _11512_/B sky130_fd_sc_hd__or2_1
XFILLER_69_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08948_ _08952_/A _08952_/B VGND VGND VPWR VPWR _08948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08879_ _08878_/Y _08866_/X _08878_/Y _08866_/X VGND VGND VPWR VPWR _08982_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10910_ _12049_/A _10910_/B VGND VGND VPWR VPWR _10910_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11890_ _11836_/A _11836_/B _11836_/Y VGND VGND VPWR VPWR _11890_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10841_ _10792_/X _10840_/Y _10792_/X _10840_/Y VGND VGND VPWR VPWR _10938_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10772_ _14563_/A _10772_/B VGND VGND VPWR VPWR _10772_/X sky130_fd_sc_hd__or2_1
XFILLER_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13560_ _13560_/A VGND VGND VPWR VPWR _13560_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12511_ _12511_/A _12511_/B VGND VGND VPWR VPWR _12511_/Y sky130_fd_sc_hd__nand2_1
X_13491_ _11516_/Y _12275_/A _11333_/Y _13490_/X VGND VGND VPWR VPWR _13491_/X sky130_fd_sc_hd__o22a_1
XFILLER_13_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15230_ _15175_/Y _15229_/Y _15175_/Y _15229_/Y VGND VGND VPWR VPWR _15285_/B sky130_fd_sc_hd__a2bb2o_1
X_12442_ _12442_/A _12442_/B VGND VGND VPWR VPWR _12442_/X sky130_fd_sc_hd__and2_1
XFILLER_40_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12373_ _12371_/A _12371_/B _12371_/X _12372_/Y VGND VGND VPWR VPWR _12437_/B sky130_fd_sc_hd__a22o_1
X_15161_ _15161_/A VGND VGND VPWR VPWR _15161_/Y sky130_fd_sc_hd__inv_2
X_14112_ _14107_/Y _14110_/Y _14111_/Y VGND VGND VPWR VPWR _14112_/X sky130_fd_sc_hd__o21a_1
X_15092_ _15075_/A _15075_/B _15075_/Y _15091_/X VGND VGND VPWR VPWR _15092_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11324_ _11324_/A VGND VGND VPWR VPWR _11324_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14043_ _14047_/A VGND VGND VPWR VPWR _14815_/A sky130_fd_sc_hd__buf_1
X_11255_ _13344_/A _11238_/B _11238_/Y _11254_/X VGND VGND VPWR VPWR _11255_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_134_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10206_ _10206_/A VGND VGND VPWR VPWR _11724_/A sky130_fd_sc_hd__clkinvlp_2
X_11186_ _11186_/A _11094_/X VGND VGND VPWR VPWR _11186_/X sky130_fd_sc_hd__or2b_1
XFILLER_79_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15994_ _15971_/X _15993_/Y _15971_/X _15993_/Y VGND VGND VPWR VPWR _16055_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10137_ _10139_/A VGND VGND VPWR VPWR _10238_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_94_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14945_ _14837_/X _14944_/Y _14844_/Y VGND VGND VPWR VPWR _14945_/X sky130_fd_sc_hd__o21a_1
X_10068_ _10067_/A _10067_/B _09971_/A _10067_/X VGND VGND VPWR VPWR _10071_/A sky130_fd_sc_hd__a22o_1
XFILLER_48_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14876_ _14876_/A VGND VGND VPWR VPWR _15544_/A sky130_fd_sc_hd__buf_1
XFILLER_90_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13827_ _14634_/A _13841_/B VGND VGND VPWR VPWR _13827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13758_ _13758_/A _13758_/B VGND VGND VPWR VPWR _13758_/X sky130_fd_sc_hd__or2_1
X_12709_ _13478_/A _12708_/X _10289_/X VGND VGND VPWR VPWR _12709_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13689_ _13675_/Y _13687_/X _13688_/Y VGND VGND VPWR VPWR _13689_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15428_ _15426_/X _15427_/Y _15426_/X _15427_/Y VGND VGND VPWR VPWR _15428_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15359_ _15420_/A _15420_/B VGND VGND VPWR VPWR _15359_/X sky130_fd_sc_hd__and2_1
XFILLER_116_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09920_ _09918_/A _09918_/B _09919_/Y VGND VGND VPWR VPWR _09921_/B sky130_fd_sc_hd__o21ai_1
XFILLER_132_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09851_ _09848_/X _09851_/B VGND VGND VPWR VPWR _09853_/B sky130_fd_sc_hd__nand2b_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08802_ _09248_/B VGND VGND VPWR VPWR _10128_/A sky130_fd_sc_hd__buf_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09782_/A _09782_/B VGND VGND VPWR VPWR _09782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08733_ _08733_/A VGND VGND VPWR VPWR _08733_/Y sky130_fd_sc_hd__inv_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08664_ _08665_/A VGND VGND VPWR VPWR _08664_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08595_ _08715_/B VGND VGND VPWR VPWR _08597_/A sky130_fd_sc_hd__buf_1
XFILLER_81_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09216_ _09216_/A VGND VGND VPWR VPWR _09216_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09147_ _08770_/A _09015_/X _08543_/B VGND VGND VPWR VPWR _09147_/X sky130_fd_sc_hd__o21ba_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09078_ _10011_/B _09078_/B VGND VGND VPWR VPWR _09165_/B sky130_fd_sc_hd__or2_1
XFILLER_123_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11040_ _10915_/X _11039_/X _10915_/X _11039_/X VGND VGND VPWR VPWR _11084_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12991_ _14488_/A _13019_/B VGND VGND VPWR VPWR _13080_/A sky130_fd_sc_hd__and2_1
XFILLER_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14730_ _14730_/A _14730_/B VGND VGND VPWR VPWR _14730_/X sky130_fd_sc_hd__or2_1
XFILLER_84_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11942_ _11942_/A _11978_/B VGND VGND VPWR VPWR _11942_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14661_ _15347_/A _14661_/B VGND VGND VPWR VPWR _14661_/Y sky130_fd_sc_hd__nand2_1
X_11873_ _11910_/A _11910_/B VGND VGND VPWR VPWR _11873_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16400_ _16407_/D VGND VGND VPWR VPWR _16400_/Y sky130_fd_sc_hd__inv_2
X_14592_ _14531_/A _14531_/B _14524_/X _14531_/Y VGND VGND VPWR VPWR _14592_/X sky130_fd_sc_hd__o2bb2a_1
X_13612_ _10421_/B _11792_/Y _10424_/B _11794_/B VGND VGND VPWR VPWR _14429_/B sky130_fd_sc_hd__o22a_1
XFILLER_60_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10824_ _12084_/A _10966_/B VGND VGND VPWR VPWR _10824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16331_ _16293_/Y _16329_/X _16330_/Y VGND VGND VPWR VPWR _16331_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13543_ _13457_/A _13494_/B _13494_/X _13542_/X VGND VGND VPWR VPWR _13543_/X sky130_fd_sc_hd__o22a_1
XFILLER_13_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10755_ _13676_/A _10631_/B _10631_/Y VGND VGND VPWR VPWR _10755_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16262_ _16262_/A _16262_/B VGND VGND VPWR VPWR _16262_/Y sky130_fd_sc_hd__nand2_1
X_13474_ _14334_/A VGND VGND VPWR VPWR _14308_/A sky130_fd_sc_hd__clkbuf_2
X_10686_ _10685_/A _10684_/Y _10685_/Y _10684_/A _10976_/A VGND VGND VPWR VPWR _10814_/B
+ sky130_fd_sc_hd__a221o_1
X_16193_ _16260_/B VGND VGND VPWR VPWR _16326_/A sky130_fd_sc_hd__buf_6
X_15213_ _15146_/A _15146_/B _15146_/Y VGND VGND VPWR VPWR _15213_/Y sky130_fd_sc_hd__o21ai_1
X_12425_ _12425_/A VGND VGND VPWR VPWR _12425_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12356_ _12305_/A _12305_/B _12305_/Y _12519_/A VGND VGND VPWR VPWR _12511_/A sky130_fd_sc_hd__a2bb2o_1
X_15144_ _15144_/A _15087_/X VGND VGND VPWR VPWR _15144_/X sky130_fd_sc_hd__or2b_1
XFILLER_126_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11307_ _13503_/A _11306_/B _11306_/X _11131_/X VGND VGND VPWR VPWR _11307_/X sky130_fd_sc_hd__o22a_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12287_ _13792_/A _12364_/B _12286_/Y VGND VGND VPWR VPWR _12287_/Y sky130_fd_sc_hd__o21ai_1
X_15075_ _15075_/A _15075_/B VGND VGND VPWR VPWR _15075_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11238_ _14038_/A _11238_/B VGND VGND VPWR VPWR _11238_/Y sky130_fd_sc_hd__nand2_1
X_14026_ _13946_/X _14025_/Y _13946_/X _14025_/Y VGND VGND VPWR VPWR _14027_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11169_ _11291_/A _11168_/Y _11291_/A _11168_/Y VGND VGND VPWR VPWR _11170_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15977_ _15984_/A _15984_/B _15976_/Y VGND VGND VPWR VPWR _15977_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14928_ _15552_/A _14928_/B VGND VGND VPWR VPWR _14928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14859_ _14859_/A _14858_/X VGND VGND VPWR VPWR _14859_/X sky130_fd_sc_hd__or2b_1
XFILLER_63_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08380_ _08380_/A VGND VGND VPWR VPWR _08401_/A sky130_fd_sc_hd__inv_2
XFILLER_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09001_ _08880_/X _09001_/B VGND VGND VPWR VPWR _09001_/X sky130_fd_sc_hd__and2b_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09903_ _09903_/A _09903_/B VGND VGND VPWR VPWR _10657_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09834_ _09834_/A VGND VGND VPWR VPWR _09834_/Y sky130_fd_sc_hd__inv_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09765_ _10049_/A VGND VGND VPWR VPWR _10079_/A sky130_fd_sc_hd__clkbuf_2
X_08716_ _08716_/A _08716_/B VGND VGND VPWR VPWR _08716_/X sky130_fd_sc_hd__or2_1
X_09696_ _09696_/A _09696_/B VGND VGND VPWR VPWR _09728_/B sky130_fd_sc_hd__or2_1
Xrebuffer30 _08662_/A VGND VGND VPWR VPWR _08380_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer41 _08368_/X VGND VGND VPWR VPWR _08414_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer52 _08398_/A VGND VGND VPWR VPWR _09232_/B sky130_fd_sc_hd__dlygate4sd1_1
X_08647_ _08647_/A VGND VGND VPWR VPWR _10110_/B sky130_fd_sc_hd__inv_2
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08578_ _09209_/A VGND VGND VPWR VPWR _10013_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10540_ _11848_/A _10540_/B VGND VGND VPWR VPWR _10540_/X sky130_fd_sc_hd__and2_1
XFILLER_50_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10471_ _10471_/A VGND VGND VPWR VPWR _10984_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12210_ _12152_/X _12209_/X _12152_/X _12209_/X VGND VGND VPWR VPWR _12211_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13190_ _13190_/A _13190_/B VGND VGND VPWR VPWR _13190_/Y sky130_fd_sc_hd__nand2_1
X_12141_ _12141_/A _12141_/B VGND VGND VPWR VPWR _12141_/X sky130_fd_sc_hd__or2_1
XFILLER_89_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12072_ _12070_/Y _12071_/Y _12010_/Y VGND VGND VPWR VPWR _12163_/A sky130_fd_sc_hd__o21ai_2
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15900_ _15900_/A _15900_/B VGND VGND VPWR VPWR _15900_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11023_ _11023_/A VGND VGND VPWR VPWR _13551_/A sky130_fd_sc_hd__buf_1
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15831_ _16238_/A VGND VGND VPWR VPWR _15832_/A sky130_fd_sc_hd__buf_6
XFILLER_66_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15762_ _15766_/A _15762_/B VGND VGND VPWR VPWR _16096_/A sky130_fd_sc_hd__or2_1
X_12974_ _12939_/X _12973_/Y _12939_/X _12973_/Y VGND VGND VPWR VPWR _13027_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14713_ _14724_/A _14724_/B VGND VGND VPWR VPWR _14807_/A sky130_fd_sc_hd__nor2_1
X_11925_ _11925_/A VGND VGND VPWR VPWR _11994_/B sky130_fd_sc_hd__inv_2
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15693_ _16053_/A VGND VGND VPWR VPWR _15693_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14644_ _14643_/A _14643_/B _11067_/B _14643_/Y VGND VGND VPWR VPWR _14644_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11856_ _11855_/A _11855_/B _11855_/X _11813_/B VGND VGND VPWR VPWR _11921_/B sky130_fd_sc_hd__a22o_1
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14575_ _14575_/A _14575_/B VGND VGND VPWR VPWR _14575_/Y sky130_fd_sc_hd__nand2_1
X_11787_ _11787_/A _11787_/B VGND VGND VPWR VPWR _11787_/X sky130_fd_sc_hd__or2_1
XFILLER_32_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10807_ _10807_/A VGND VGND VPWR VPWR _10807_/Y sky130_fd_sc_hd__inv_2
X_16314_ _16248_/Y _16313_/Y _16248_/Y _16313_/Y VGND VGND VPWR VPWR _16316_/B sky130_fd_sc_hd__o2bb2a_1
X_10738_ _11970_/A VGND VGND VPWR VPWR _13083_/A sky130_fd_sc_hd__buf_1
X_13526_ _10326_/X _13481_/X _10326_/X _13481_/X VGND VGND VPWR VPWR _13527_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16245_ _16245_/A _15785_/X VGND VGND VPWR VPWR _16246_/A sky130_fd_sc_hd__or2b_1
X_13457_ _13457_/A _13457_/B VGND VGND VPWR VPWR _13457_/Y sky130_fd_sc_hd__nor2_1
X_12408_ _14005_/A _12407_/B _12407_/Y VGND VGND VPWR VPWR _12408_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10669_ _09984_/A _09984_/B _09984_/Y VGND VGND VPWR VPWR _10670_/A sky130_fd_sc_hd__o21ai_1
XFILLER_126_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16176_ _16192_/A _16176_/B VGND VGND VPWR VPWR _16264_/B sky130_fd_sc_hd__or2_1
XFILLER_114_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13388_ _13363_/X _13387_/X _13363_/X _13387_/X VGND VGND VPWR VPWR _13439_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12339_ _14028_/A _12223_/B _12223_/Y VGND VGND VPWR VPWR _12339_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15127_ _15093_/X _15126_/Y _15093_/X _15126_/Y VGND VGND VPWR VPWR _15128_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15058_ _15058_/A _15044_/X VGND VGND VPWR VPWR _15058_/X sky130_fd_sc_hd__or2b_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14009_ _15416_/A _13957_/B _13957_/Y VGND VGND VPWR VPWR _14009_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09550_ _09613_/A _09548_/X _09613_/B VGND VGND VPWR VPWR _09550_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09481_ _08757_/A _09477_/X _08757_/A _09477_/X VGND VGND VPWR VPWR _09482_/B sky130_fd_sc_hd__o2bb2a_1
X_08501_ _08501_/A VGND VGND VPWR VPWR _08501_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_64_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08432_ _08713_/A VGND VGND VPWR VPWR _09323_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08363_ input27/X _08363_/B VGND VGND VPWR VPWR _08364_/B sky130_fd_sc_hd__nor2_1
X_08294_ _08311_/A input21/X _08312_/A _08314_/A VGND VGND VPWR VPWR _08309_/A sky130_fd_sc_hd__o22a_1
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09817_ _09817_/A _09817_/B _09826_/B VGND VGND VPWR VPWR _09818_/B sky130_fd_sc_hd__or3_1
XFILLER_100_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09748_ _09748_/A VGND VGND VPWR VPWR _10034_/A sky130_fd_sc_hd__inv_2
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A VGND VGND VPWR VPWR _11710_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09679_ _09679_/A1 _09681_/B _09799_/B VGND VGND VPWR VPWR _09829_/B sky130_fd_sc_hd__o21ai_2
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12690_ _10826_/A _12669_/A _10826_/Y _12669_/Y VGND VGND VPWR VPWR _12691_/B sky130_fd_sc_hd__o22a_1
XFILLER_15_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _12390_/A _11641_/B VGND VGND VPWR VPWR _11641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14360_ _14377_/A _14377_/B VGND VGND VPWR VPWR _14360_/Y sky130_fd_sc_hd__nor2_1
X_11572_ _11572_/A _11572_/B VGND VGND VPWR VPWR _14148_/A sky130_fd_sc_hd__or2_1
XFILLER_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13311_ _14858_/A _13306_/B _13306_/Y VGND VGND VPWR VPWR _13311_/Y sky130_fd_sc_hd__o21ai_1
X_10523_ _11836_/A _10523_/B VGND VGND VPWR VPWR _10523_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 wbs_dat_i[10] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__buf_1
XFILLER_10_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14291_ _13447_/A _13447_/B _13447_/Y VGND VGND VPWR VPWR _14291_/X sky130_fd_sc_hd__o21a_1
X_16030_ _16030_/A _16030_/B VGND VGND VPWR VPWR _16030_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13242_ _14438_/A VGND VGND VPWR VPWR _14732_/A sky130_fd_sc_hd__buf_1
X_10454_ _10454_/A VGND VGND VPWR VPWR _10968_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13173_ _13104_/X _13172_/Y _13104_/X _13172_/Y VGND VGND VPWR VPWR _13186_/B sky130_fd_sc_hd__a2bb2o_1
X_10385_ _10251_/A _10384_/Y _10251_/Y _10384_/A _10471_/A VGND VGND VPWR VPWR _11806_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_6_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12124_ _13917_/A _12145_/B VGND VGND VPWR VPWR _12221_/A sky130_fd_sc_hd__and2_1
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12055_ _12055_/A _12055_/B VGND VGND VPWR VPWR _12055_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11006_ _11006_/A _11005_/X VGND VGND VPWR VPWR _11006_/X sky130_fd_sc_hd__or2b_1
XFILLER_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15814_ _15737_/Y _15812_/X _15813_/Y VGND VGND VPWR VPWR _15814_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15745_ _14915_/X _15744_/X _14915_/X _15744_/X VGND VGND VPWR VPWR _15746_/B sky130_fd_sc_hd__a2bb2oi_1
X_12957_ _14944_/A _12949_/B _12949_/Y VGND VGND VPWR VPWR _12957_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15676_ _15622_/Y _15674_/X _15675_/Y VGND VGND VPWR VPWR _15676_/X sky130_fd_sc_hd__o21a_1
X_11908_ _11876_/Y _11906_/Y _11907_/Y VGND VGND VPWR VPWR _11909_/A sky130_fd_sc_hd__o21ai_2
X_12888_ _14476_/A _12938_/B VGND VGND VPWR VPWR _12888_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14627_ _14579_/A _14579_/B _14579_/Y VGND VGND VPWR VPWR _14627_/Y sky130_fd_sc_hd__o21ai_1
X_11839_ _11833_/Y _11837_/X _11838_/Y VGND VGND VPWR VPWR _11839_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14558_ _14577_/A _14577_/B VGND VGND VPWR VPWR _14558_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14489_ _14464_/A _14464_/B _14464_/Y VGND VGND VPWR VPWR _14489_/Y sky130_fd_sc_hd__o21ai_1
X_13509_ _13509_/A _13509_/B VGND VGND VPWR VPWR _13509_/Y sky130_fd_sc_hd__nand2_1
X_16228_ _16228_/A VGND VGND VPWR VPWR _16228_/Y sky130_fd_sc_hd__inv_2
X_16159_ _15816_/X _16158_/X _15816_/X _16158_/X VGND VGND VPWR VPWR _16160_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08981_ _08885_/X _08979_/X _11359_/B VGND VGND VPWR VPWR _08981_/X sky130_fd_sc_hd__o21a_2
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09602_ _09552_/X _09601_/Y _09552_/X _09601_/Y VGND VGND VPWR VPWR _09656_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09533_ _09555_/A _09555_/B VGND VGND VPWR VPWR _09595_/A sky130_fd_sc_hd__nor2_1
XFILLER_71_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09464_ _10017_/A _08623_/A _09457_/Y _09463_/X VGND VGND VPWR VPWR _09464_/X sky130_fd_sc_hd__o22a_1
X_09395_ _09395_/A VGND VGND VPWR VPWR _13648_/A sky130_fd_sc_hd__buf_1
XFILLER_52_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08415_ _08415_/A1 _08348_/Y _08414_/Y _08348_/A _08419_/A VGND VGND VPWR VPWR _09221_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08346_ input29/X _08346_/B VGND VGND VPWR VPWR _08347_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08277_ input25/X VGND VGND VPWR VPWR _08278_/A sky130_fd_sc_hd__inv_2
XFILLER_20_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10170_ _10251_/A _10170_/B VGND VGND VPWR VPWR _10170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13860_ _13799_/Y _13858_/X _13859_/Y VGND VGND VPWR VPWR _13860_/X sky130_fd_sc_hd__o21a_1
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13791_ _13792_/A _13792_/B VGND VGND VPWR VPWR _13791_/X sky130_fd_sc_hd__and2_1
X_12811_ _12849_/A _12849_/B VGND VGND VPWR VPWR _12811_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15530_ _15526_/Y _15624_/A _15529_/Y VGND VGND VPWR VPWR _15534_/B sky130_fd_sc_hd__o21ai_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12776_/A _12776_/B VGND VGND VPWR VPWR _12742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15461_ _15461_/A _15461_/B VGND VGND VPWR VPWR _15461_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12673_ _12673_/A VGND VGND VPWR VPWR _12673_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _10424_/A _10421_/B _12833_/A _11720_/B VGND VGND VPWR VPWR _14412_/X sky130_fd_sc_hd__a22o_1
X_11624_ _11621_/Y _12419_/A _11520_/X _11623_/Y VGND VGND VPWR VPWR _11624_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15392_ _15392_/A _15398_/B VGND VGND VPWR VPWR _15468_/A sky130_fd_sc_hd__and2_1
XFILLER_128_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14343_ _14255_/A _14342_/Y _14255_/A _14342_/Y VGND VGND VPWR VPWR _14381_/A sky130_fd_sc_hd__a2bb2o_1
X_11555_ _12400_/A _11557_/B VGND VGND VPWR VPWR _11558_/A sky130_fd_sc_hd__and2_1
XFILLER_11_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14274_ _15857_/A _14274_/B VGND VGND VPWR VPWR _14274_/Y sky130_fd_sc_hd__nand2_1
X_11486_ _11586_/A _11486_/B VGND VGND VPWR VPWR _13206_/A sky130_fd_sc_hd__or2_2
X_10506_ _09832_/A _09832_/B _09833_/A VGND VGND VPWR VPWR _10507_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16013_ _16038_/A _16038_/B VGND VGND VPWR VPWR _16013_/Y sky130_fd_sc_hd__nor2_1
X_13225_ _14740_/A _13300_/B VGND VGND VPWR VPWR _13225_/Y sky130_fd_sc_hd__nor2_1
X_10437_ _10437_/A VGND VGND VPWR VPWR _10437_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13156_ _13198_/A _13198_/B VGND VGND VPWR VPWR _13156_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10368_ _10365_/Y _12701_/A _10299_/X _10367_/Y VGND VGND VPWR VPWR _10368_/X sky130_fd_sc_hd__o22a_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12107_ _13200_/A _12157_/B _12106_/Y VGND VGND VPWR VPWR _12107_/Y sky130_fd_sc_hd__o21ai_1
X_13087_ _15261_/A _13107_/B VGND VGND VPWR VPWR _13087_/Y sky130_fd_sc_hd__nor2_1
X_10299_ _10296_/A _10325_/B _10295_/X _10298_/Y VGND VGND VPWR VPWR _10299_/X sky130_fd_sc_hd__o22a_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12038_ _11967_/X _12037_/Y _11967_/X _12037_/Y VGND VGND VPWR VPWR _12053_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_120_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13989_ _14956_/A _13988_/B _13988_/Y VGND VGND VPWR VPWR _13989_/X sky130_fd_sc_hd__a21o_1
X_15728_ _15728_/A _15728_/B VGND VGND VPWR VPWR _16114_/A sky130_fd_sc_hd__nor2_1
XFILLER_46_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15659_ _12611_/A _15658_/A _12611_/Y _15658_/Y _15655_/B VGND VGND VPWR VPWR _16027_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09180_ _09431_/A _09180_/B VGND VGND VPWR VPWR _09180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08964_ _08963_/Y _08859_/X _08963_/Y _08859_/X VGND VGND VPWR VPWR _08968_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_130_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08895_ _08894_/Y _08863_/X _08894_/Y _08863_/X VGND VGND VPWR VPWR _08976_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09516_ _09484_/A _09484_/B _09484_/Y _09515_/X VGND VGND VPWR VPWR _09516_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _12065_/A VGND VGND VPWR VPWR _10924_/A sky130_fd_sc_hd__inv_2
XFILLER_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09378_ _09354_/X _09377_/X _09354_/X _09377_/X VGND VGND VPWR VPWR _09379_/A sky130_fd_sc_hd__a2bb2o_1
X_08329_ _08329_/A VGND VGND VPWR VPWR _08329_/Y sky130_fd_sc_hd__inv_2
X_11340_ _13780_/A _11500_/B VGND VGND VPWR VPWR _11340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13010_ _14504_/A _13010_/B VGND VGND VPWR VPWR _13010_/Y sky130_fd_sc_hd__nor2_1
X_11271_ _11271_/A _11271_/B VGND VGND VPWR VPWR _11271_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10222_ _10222_/A VGND VGND VPWR VPWR _10222_/Y sky130_fd_sc_hd__inv_2
X_10153_ _10155_/A VGND VGND VPWR VPWR _10242_/B sky130_fd_sc_hd__buf_1
XFILLER_121_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14961_ _14971_/A _14971_/B VGND VGND VPWR VPWR _14961_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10084_ _10043_/X _10082_/X _11142_/B VGND VGND VPWR VPWR _10084_/X sky130_fd_sc_hd__o21a_1
X_14892_ _15529_/A _14912_/B VGND VGND VPWR VPWR _14892_/Y sky130_fd_sc_hd__nor2_1
X_13912_ _15408_/A _13949_/B VGND VGND VPWR VPWR _13912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13843_ _14630_/A _13843_/B VGND VGND VPWR VPWR _13843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15513_ _15470_/A _15470_/B _15470_/Y VGND VGND VPWR VPWR _15513_/Y sky130_fd_sc_hd__o21ai_1
X_13774_ _13774_/A _13774_/B VGND VGND VPWR VPWR _13800_/B sky130_fd_sc_hd__or2_1
X_10986_ _12174_/A VGND VGND VPWR VPWR _12689_/A sky130_fd_sc_hd__buf_1
XFILLER_16_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12725_ _12683_/A _12683_/B _12683_/Y VGND VGND VPWR VPWR _12725_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15444_ _15444_/A _15414_/X VGND VGND VPWR VPWR _15444_/X sky130_fd_sc_hd__or2b_1
X_12656_ _12864_/A VGND VGND VPWR VPWR _15171_/A sky130_fd_sc_hd__buf_1
XFILLER_31_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12587_ _12587_/A _11431_/X VGND VGND VPWR VPWR _12588_/A sky130_fd_sc_hd__or2b_1
X_15375_ _15375_/A _15341_/X VGND VGND VPWR VPWR _15375_/X sky130_fd_sc_hd__or2b_1
X_11607_ _11607_/A _11607_/B VGND VGND VPWR VPWR _12426_/A sky130_fd_sc_hd__or2_1
XFILLER_128_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14326_ _14111_/A _13435_/B _13435_/Y VGND VGND VPWR VPWR _14326_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11538_ _11623_/A _12419_/A VGND VGND VPWR VPWR _11538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14257_ _14221_/Y _14255_/Y _14256_/Y VGND VGND VPWR VPWR _14258_/A sky130_fd_sc_hd__o21ai_1
X_11469_ _09430_/A _09185_/B _09185_/Y VGND VGND VPWR VPWR _11470_/A sky130_fd_sc_hd__o21ai_1
X_14188_ _14206_/A _14188_/B VGND VGND VPWR VPWR _15860_/A sky130_fd_sc_hd__or2_1
X_13208_ _13140_/X _13207_/X _13140_/X _13207_/X VGND VGND VPWR VPWR _13451_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_98_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13139_ _13139_/A _13139_/B VGND VGND VPWR VPWR _13139_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08680_ _08679_/A _08679_/B _08678_/Y _08679_/X VGND VGND VPWR VPWR _08680_/X sky130_fd_sc_hd__o22a_1
XFILLER_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09301_ _09300_/A _08946_/Y _09300_/Y _08946_/A VGND VGND VPWR VPWR _10235_/A sky130_fd_sc_hd__o22a_1
XFILLER_34_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09232_ _09232_/A _09232_/B VGND VGND VPWR VPWR _09400_/A sky130_fd_sc_hd__or2_1
X_09163_ _08757_/Y _09160_/A _08757_/A _09160_/Y VGND VGND VPWR VPWR _10009_/B sky130_fd_sc_hd__o22a_1
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09094_ _09705_/A VGND VGND VPWR VPWR _09415_/A sky130_fd_sc_hd__buf_1
XFILLER_134_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09996_ _09965_/X _11309_/A _11308_/B VGND VGND VPWR VPWR _11513_/A sky130_fd_sc_hd__o21a_1
XFILLER_97_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08947_ _08946_/Y _08857_/X _08946_/Y _08857_/X VGND VGND VPWR VPWR _08952_/B sky130_fd_sc_hd__o2bb2a_1
X_08878_ _08770_/A _10132_/A _08770_/Y VGND VGND VPWR VPWR _08878_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10840_ _13640_/A _10946_/B _10839_/Y VGND VGND VPWR VPWR _10840_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10771_ _11966_/A VGND VGND VPWR VPWR _14563_/A sky130_fd_sc_hd__buf_1
X_12510_ _13445_/A _12302_/B _12302_/Y VGND VGND VPWR VPWR _12511_/B sky130_fd_sc_hd__o21a_1
XFILLER_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13490_ _11311_/Y _12181_/A _11157_/Y _13489_/X VGND VGND VPWR VPWR _13490_/X sky130_fd_sc_hd__o22a_1
X_12441_ _13462_/A _12441_/B VGND VGND VPWR VPWR _12441_/X sky130_fd_sc_hd__and2_1
XFILLER_12_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12372_ _12372_/A VGND VGND VPWR VPWR _12372_/Y sky130_fd_sc_hd__inv_2
X_15160_ _12381_/X _15101_/X _12383_/B VGND VGND VPWR VPWR _15161_/A sky130_fd_sc_hd__o21ai_2
XFILLER_4_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14111_ _14111_/A _14111_/B VGND VGND VPWR VPWR _14111_/Y sky130_fd_sc_hd__nand2_1
X_15091_ _15078_/A _15078_/B _15078_/Y _15090_/X VGND VGND VPWR VPWR _15091_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11323_ _11323_/A VGND VGND VPWR VPWR _11323_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14042_ _14042_/A _14042_/B VGND VGND VPWR VPWR _14042_/Y sky130_fd_sc_hd__nor2_1
X_11254_ _13348_/A _11244_/B _11244_/Y _11253_/X VGND VGND VPWR VPWR _11254_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10205_ _10346_/B _10902_/B VGND VGND VPWR VPWR _10206_/A sky130_fd_sc_hd__or2_1
X_11185_ _14059_/A VGND VGND VPWR VPWR _15446_/A sky130_fd_sc_hd__buf_1
XFILLER_69_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15993_ _15915_/X _15993_/B VGND VGND VPWR VPWR _15993_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10136_ _10120_/A _10120_/B _10120_/X VGND VGND VPWR VPWR _10139_/A sky130_fd_sc_hd__a21bo_1
XFILLER_121_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14944_ _14944_/A _14944_/B VGND VGND VPWR VPWR _14944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10067_ _10067_/A _10067_/B VGND VGND VPWR VPWR _10067_/X sky130_fd_sc_hd__or2_1
XFILLER_48_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14875_ _15546_/A _14922_/B VGND VGND VPWR VPWR _14875_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13826_ _13757_/X _13825_/X _13757_/X _13825_/X VGND VGND VPWR VPWR _13841_/B sky130_fd_sc_hd__a2bb2o_1
X_13757_ _13749_/Y _13755_/X _13756_/Y VGND VGND VPWR VPWR _13757_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10969_ _10046_/X _10969_/B VGND VGND VPWR VPWR _10969_/X sky130_fd_sc_hd__and2b_1
X_12708_ _10284_/Y _10350_/B _12708_/B1 _10349_/A VGND VGND VPWR VPWR _12708_/X sky130_fd_sc_hd__o22a_1
X_13688_ _14496_/A _13688_/B VGND VGND VPWR VPWR _13688_/Y sky130_fd_sc_hd__nand2_1
X_15427_ _12431_/A _15163_/B _15163_/Y _15165_/Y VGND VGND VPWR VPWR _15427_/Y sky130_fd_sc_hd__o2bb2ai_1
X_12639_ _14283_/A _12637_/X _12638_/X VGND VGND VPWR VPWR _12639_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15358_ _15352_/X _15357_/Y _15352_/X _15357_/Y VGND VGND VPWR VPWR _15420_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14309_ _15857_/A _14274_/B _14274_/Y VGND VGND VPWR VPWR _14309_/Y sky130_fd_sc_hd__o21ai_1
X_15289_ _15289_/A _15289_/B VGND VGND VPWR VPWR _15289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09850_ _09848_/A _09848_/B _09849_/Y VGND VGND VPWR VPWR _09851_/B sky130_fd_sc_hd__o21ai_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08801_ _08801_/A VGND VGND VPWR VPWR _09248_/B sky130_fd_sc_hd__inv_2
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09782_/A _09782_/B VGND VGND VPWR VPWR _09781_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08732_ _08713_/A _08713_/B _08713_/X _08731_/Y VGND VGND VPWR VPWR _08733_/A sky130_fd_sc_hd__a22o_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08663_ _09677_/A _08663_/B VGND VGND VPWR VPWR _08665_/A sky130_fd_sc_hd__or2_1
XFILLER_54_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08594_ _09455_/B VGND VGND VPWR VPWR _08715_/B sky130_fd_sc_hd__inv_2
XFILLER_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09215_ _09551_/A _09728_/A VGND VGND VPWR VPWR _09216_/A sky130_fd_sc_hd__or2_1
XFILLER_14_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09146_ _09146_/A VGND VGND VPWR VPWR _09146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09077_ _10012_/B _09077_/B VGND VGND VPWR VPWR _09078_/B sky130_fd_sc_hd__or2_1
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09979_ _09970_/Y _09977_/Y _09978_/Y VGND VGND VPWR VPWR _09981_/B sky130_fd_sc_hd__o21ai_1
XFILLER_76_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12990_ _12931_/X _12989_/Y _12931_/X _12989_/Y VGND VGND VPWR VPWR _13019_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11941_ _11981_/A _11940_/Y _11981_/A _11940_/Y VGND VGND VPWR VPWR _11978_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14660_ _14613_/Y _14658_/X _14659_/Y VGND VGND VPWR VPWR _14660_/X sky130_fd_sc_hd__o21a_1
X_11872_ _11847_/X _11871_/Y _11847_/X _11871_/Y VGND VGND VPWR VPWR _11910_/B sky130_fd_sc_hd__a2bb2o_1
X_13611_ _13611_/A VGND VGND VPWR VPWR _13611_/Y sky130_fd_sc_hd__inv_2
X_14591_ _14591_/A VGND VGND VPWR VPWR _15187_/A sky130_fd_sc_hd__buf_1
X_10823_ _10822_/A _10821_/Y _10822_/Y _10821_/A _10976_/A VGND VGND VPWR VPWR _10966_/B
+ sky130_fd_sc_hd__a221o_1
X_16330_ _16330_/A _16330_/B VGND VGND VPWR VPWR _16330_/Y sky130_fd_sc_hd__nand2_1
X_13542_ _15104_/A _13497_/B _13497_/Y _13541_/X VGND VGND VPWR VPWR _13542_/X sky130_fd_sc_hd__a2bb2o_1
X_10754_ _11895_/A VGND VGND VPWR VPWR _13676_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16261_ _16194_/Y _16259_/X _16260_/Y VGND VGND VPWR VPWR _16261_/X sky130_fd_sc_hd__o21a_1
X_13473_ _14352_/A VGND VGND VPWR VPWR _14334_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10685_ _10685_/A VGND VGND VPWR VPWR _10685_/Y sky130_fd_sc_hd__inv_2
X_16192_ _16192_/A _16192_/B VGND VGND VPWR VPWR _16260_/B sky130_fd_sc_hd__or2_1
X_15212_ _15212_/A _15212_/B VGND VGND VPWR VPWR _15212_/X sky130_fd_sc_hd__or2_1
X_12424_ _12435_/B VGND VGND VPWR VPWR _12424_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12355_ _12308_/A _12308_/B _12308_/Y _12527_/A VGND VGND VPWR VPWR _12519_/A sky130_fd_sc_hd__a2bb2o_1
X_15143_ _15143_/A _15143_/B VGND VGND VPWR VPWR _15143_/Y sky130_fd_sc_hd__nand2_1
X_11306_ _12172_/A _11306_/B VGND VGND VPWR VPWR _11306_/X sky130_fd_sc_hd__and2_1
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12286_ _12364_/A _12364_/B VGND VGND VPWR VPWR _12286_/Y sky130_fd_sc_hd__nand2_1
X_15074_ _15033_/X _15073_/X _15033_/X _15073_/X VGND VGND VPWR VPWR _15075_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11237_ _11079_/X _11236_/X _11079_/X _11236_/X VGND VGND VPWR VPWR _11238_/B sky130_fd_sc_hd__a2bb2o_1
X_14025_ _15406_/A _13947_/B _13947_/Y VGND VGND VPWR VPWR _14025_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11168_ _13719_/A _11290_/B _11167_/Y VGND VGND VPWR VPWR _11168_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10119_ _10119_/A _10119_/B VGND VGND VPWR VPWR _10120_/A sky130_fd_sc_hd__or2_1
X_15976_ _15984_/A _15984_/B VGND VGND VPWR VPWR _15976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11099_ _11304_/A VGND VGND VPWR VPWR _12261_/A sky130_fd_sc_hd__buf_1
XFILLER_48_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14927_ _14867_/Y _14925_/X _14926_/Y VGND VGND VPWR VPWR _14927_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14858_ _14858_/A _14858_/B VGND VGND VPWR VPWR _14858_/X sky130_fd_sc_hd__or2_1
XFILLER_63_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13809_ _13809_/A _13768_/X VGND VGND VPWR VPWR _13809_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14789_ _14733_/X _14788_/X _14733_/X _14788_/X VGND VGND VPWR VPWR _14790_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16459_ _16357_/A _16459_/D VGND VGND VPWR VPWR _16459_/Q sky130_fd_sc_hd__dfxtp_1
X_09000_ _11393_/A VGND VGND VPWR VPWR _11572_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09902_ _09903_/A _09903_/B VGND VGND VPWR VPWR _10657_/B sky130_fd_sc_hd__and2_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _09833_/A VGND VGND VPWR VPWR _09833_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09733_/A _09733_/B _09736_/A VGND VGND VPWR VPWR _10049_/A sky130_fd_sc_hd__a21bo_1
XFILLER_27_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08715_ _08715_/A _08715_/B VGND VGND VPWR VPWR _08715_/X sky130_fd_sc_hd__or2_1
X_09695_ _09695_/A _09695_/B VGND VGND VPWR VPWR _09698_/A sky130_fd_sc_hd__or2_1
Xrebuffer20 rebuffer21/X VGND VGND VPWR VPWR rebuffer20/X sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08646_ _08645_/X _08407_/Y _08645_/X _08407_/Y VGND VGND VPWR VPWR _08647_/A sky130_fd_sc_hd__o2bb2a_1
Xrebuffer53 rebuffer57/X VGND VGND VPWR VPWR _09005_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer42 _10189_/X VGND VGND VPWR VPWR _11148_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer31 _10173_/A VGND VGND VPWR VPWR _10304_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _09454_/B VGND VGND VPWR VPWR _09553_/A sky130_fd_sc_hd__buf_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10470_ _10470_/A VGND VGND VPWR VPWR _10470_/Y sky130_fd_sc_hd__clkinvlp_2
X_09129_ _09553_/B _09035_/B _09036_/B VGND VGND VPWR VPWR _09130_/A sky130_fd_sc_hd__a21bo_1
X_12140_ _12230_/A _12138_/X _12139_/X VGND VGND VPWR VPWR _12140_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12071_ _12071_/A VGND VGND VPWR VPWR _12071_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11022_ _13905_/A _11090_/B VGND VGND VPWR VPWR _11204_/A sky130_fd_sc_hd__and2_1
X_15830_ _14406_/Y _15829_/X _14406_/Y _15829_/X VGND VGND VPWR VPWR _16238_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_106_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15761_ _14909_/X _15760_/X _14909_/X _15760_/X VGND VGND VPWR VPWR _15762_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12973_ _14531_/A _12940_/B _12940_/Y VGND VGND VPWR VPWR _12973_/Y sky130_fd_sc_hd__o21ai_1
X_15692_ _15700_/A _15692_/B VGND VGND VPWR VPWR _16053_/A sky130_fd_sc_hd__or2_1
X_14712_ _14646_/Y _14711_/Y _14646_/Y _14711_/Y VGND VGND VPWR VPWR _14724_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11924_ _10561_/A _11859_/A _10677_/B _11923_/Y VGND VGND VPWR VPWR _11925_/A sky130_fd_sc_hd__o22a_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14643_ _14643_/A _14643_/B VGND VGND VPWR VPWR _14643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11855_ _11855_/A _11855_/B VGND VGND VPWR VPWR _11855_/X sky130_fd_sc_hd__or2_1
XFILLER_33_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14574_ _14566_/Y _14572_/X _14573_/Y VGND VGND VPWR VPWR _14574_/X sky130_fd_sc_hd__o21a_1
X_11786_ _11787_/A _11787_/B VGND VGND VPWR VPWR _11788_/A sky130_fd_sc_hd__and2_1
X_10806_ _09987_/A _09987_/B _09987_/Y VGND VGND VPWR VPWR _10807_/A sky130_fd_sc_hd__o21ai_1
XFILLER_32_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16313_ _16249_/A _16316_/A _16249_/Y VGND VGND VPWR VPWR _16313_/Y sky130_fd_sc_hd__o21ai_1
X_13525_ _13527_/A VGND VGND VPWR VPWR _15030_/A sky130_fd_sc_hd__buf_1
XFILLER_41_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10737_ _10735_/A _10736_/A _10735_/Y _10736_/Y _09672_/A VGND VGND VPWR VPWR _11970_/A
+ sky130_fd_sc_hd__a221o_2
X_16244_ _16244_/A VGND VGND VPWR VPWR _16457_/S sky130_fd_sc_hd__clkbuf_2
X_13456_ _13130_/X _13455_/X _13130_/X _13455_/X VGND VGND VPWR VPWR _13456_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12407_ _14005_/A _12407_/B VGND VGND VPWR VPWR _12407_/Y sky130_fd_sc_hd__nand2_1
X_10668_ _13515_/A _10667_/B _10667_/X _10547_/X VGND VGND VPWR VPWR _10668_/X sky130_fd_sc_hd__o22a_1
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16175_ _15812_/X _16174_/X _15812_/X _16174_/X VGND VGND VPWR VPWR _16176_/B sky130_fd_sc_hd__a2bb2o_1
X_13387_ _13387_/A _13364_/X VGND VGND VPWR VPWR _13387_/X sky130_fd_sc_hd__or2b_1
X_10599_ _09963_/Y _10598_/A _09963_/A _10598_/Y _09797_/A VGND VGND VPWR VPWR _11882_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_126_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12338_ _13395_/A _12341_/B VGND VGND VPWR VPWR _12338_/Y sky130_fd_sc_hd__nor2_1
X_15126_ _15069_/A _15069_/B _15069_/Y VGND VGND VPWR VPWR _15126_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15057_ _15057_/A _15057_/B VGND VGND VPWR VPWR _15057_/Y sky130_fd_sc_hd__nand2_1
X_12269_ _12687_/A _12268_/B _12268_/X _12181_/B VGND VGND VPWR VPWR _12376_/B sky130_fd_sc_hd__a22o_1
X_14008_ _14008_/A _14063_/B VGND VGND VPWR VPWR _14008_/X sky130_fd_sc_hd__and2_1
XFILLER_110_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15959_ _15930_/X _15957_/X _16008_/B VGND VGND VPWR VPWR _15959_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08500_ _08589_/A VGND VGND VPWR VPWR _08701_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09480_ _08749_/A _09520_/S _08749_/A _09520_/S VGND VGND VPWR VPWR _09518_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08431_ _09209_/A VGND VGND VPWR VPWR _08713_/A sky130_fd_sc_hd__inv_2
XFILLER_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08362_ _08275_/A input10/X _08387_/B _08361_/Y VGND VGND VPWR VPWR _08366_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08293_ _08316_/A input20/X _08317_/A _08319_/A VGND VGND VPWR VPWR _08314_/A sky130_fd_sc_hd__o22a_1
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09816_ _09809_/X _08839_/Y _09809_/X _08839_/Y VGND VGND VPWR VPWR _09818_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09747_ _09791_/A _09791_/B _09791_/A _09791_/B VGND VGND VPWR VPWR _09748_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09678_ _09707_/B _09680_/A VGND VGND VPWR VPWR _09799_/B sky130_fd_sc_hd__or2_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08629_ _09458_/B VGND VGND VPWR VPWR _09538_/A sky130_fd_sc_hd__buf_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A _11639_/X VGND VGND VPWR VPWR _11640_/X sky130_fd_sc_hd__or2b_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11571_ _08985_/X _11570_/X _08985_/X _11570_/X VGND VGND VPWR VPWR _11572_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_128_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13310_ _14067_/A _13309_/B _13309_/Y VGND VGND VPWR VPWR _13310_/X sky130_fd_sc_hd__a21o_1
X_10522_ _10522_/A VGND VGND VPWR VPWR _10522_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14290_ _15982_/A _14404_/B VGND VGND VPWR VPWR _14290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13241_ _15069_/A VGND VGND VPWR VPWR _14438_/A sky130_fd_sc_hd__inv_2
X_10453_ _10452_/Y _10370_/X _10379_/Y VGND VGND VPWR VPWR _10453_/X sky130_fd_sc_hd__o21a_1
X_13172_ _15264_/A _13105_/B _13105_/Y VGND VGND VPWR VPWR _13172_/Y sky130_fd_sc_hd__o21ai_1
X_10384_ _10384_/A VGND VGND VPWR VPWR _10384_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12123_ _12056_/X _12122_/Y _12056_/X _12122_/Y VGND VGND VPWR VPWR _12145_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12054_ _12039_/Y _12052_/X _12053_/Y VGND VGND VPWR VPWR _12054_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11005_ _14409_/A _11005_/B VGND VGND VPWR VPWR _11005_/X sky130_fd_sc_hd__or2_1
X_15813_ _16112_/A _15813_/B VGND VGND VPWR VPWR _15813_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15744_ _14916_/A _14916_/B _14916_/Y VGND VGND VPWR VPWR _15744_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12956_ _13878_/A VGND VGND VPWR VPWR _14836_/A sky130_fd_sc_hd__buf_1
XFILLER_61_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15675_ _15675_/A _15675_/B VGND VGND VPWR VPWR _15675_/Y sky130_fd_sc_hd__nand2_1
X_11907_ _11907_/A _11907_/B VGND VGND VPWR VPWR _11907_/Y sky130_fd_sc_hd__nand2_1
X_12887_ _12850_/X _12886_/Y _12850_/X _12886_/Y VGND VGND VPWR VPWR _12938_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14626_/A VGND VGND VPWR VPWR _15337_/A sky130_fd_sc_hd__buf_1
X_11838_ _11838_/A _11838_/B VGND VGND VPWR VPWR _11838_/Y sky130_fd_sc_hd__nand2_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14512_/X _14556_/X _14512_/X _14556_/X VGND VGND VPWR VPWR _14577_/B sky130_fd_sc_hd__a2bb2o_1
X_11769_ _11806_/B _11768_/Y _11806_/B _11768_/Y VGND VGND VPWR VPWR _11802_/A sky130_fd_sc_hd__a2bb2o_1
X_13508_ _10833_/X _13487_/X _10833_/X _13487_/X VGND VGND VPWR VPWR _13509_/B sky130_fd_sc_hd__o2bb2a_1
X_14488_ _14488_/A VGND VGND VPWR VPWR _15202_/A sky130_fd_sc_hd__buf_1
X_16227_ _16227_/A VGND VGND VPWR VPWR _16227_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_127_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13439_ _13439_/A _13439_/B VGND VGND VPWR VPWR _13439_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16158_ _15817_/A _15817_/B _15817_/Y VGND VGND VPWR VPWR _16158_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15109_ _15099_/X _15108_/Y _15099_/X _15108_/Y VGND VGND VPWR VPWR _15110_/B sky130_fd_sc_hd__a2bb2o_1
X_16089_ _16089_/A _16089_/B VGND VGND VPWR VPWR _16089_/Y sky130_fd_sc_hd__nand2_1
X_08980_ _08980_/A _08980_/B VGND VGND VPWR VPWR _11359_/B sky130_fd_sc_hd__or2_1
XFILLER_87_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09601_ _09601_/A _09601_/B VGND VGND VPWR VPWR _09601_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09532_ _09532_/A VGND VGND VPWR VPWR _09532_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09463_ _09458_/Y _09461_/X _09462_/X VGND VGND VPWR VPWR _09463_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09394_ _11128_/A VGND VGND VPWR VPWR _09395_/A sky130_fd_sc_hd__buf_1
XFILLER_51_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08414_ _08414_/A VGND VGND VPWR VPWR _08414_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08345_ _08343_/Y _08344_/A _08343_/A _08344_/Y _08304_/A VGND VGND VPWR VPWR _09217_/B
+ sky130_fd_sc_hd__o221a_1
X_08276_ input9/X VGND VGND VPWR VPWR _08276_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12810_ _12773_/X _12809_/Y _12773_/X _12809_/Y VGND VGND VPWR VPWR _12849_/B sky130_fd_sc_hd__a2bb2o_1
X_13790_ _13863_/A _13789_/Y _13863_/A _13789_/Y VGND VGND VPWR VPWR _13792_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12715_/X _12740_/X _12715_/X _12740_/X VGND VGND VPWR VPWR _12776_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15460_ _15403_/X _15459_/X _15403_/X _15459_/X VGND VGND VPWR VPWR _15461_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _11140_/Y _12671_/Y _10978_/Y VGND VGND VPWR VPWR _12673_/A sky130_fd_sc_hd__o21ai_1
X_14411_ _14411_/A VGND VGND VPWR VPWR _15193_/A sky130_fd_sc_hd__buf_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A _12382_/A VGND VGND VPWR VPWR _11623_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15391_ _15330_/X _15390_/Y _15330_/X _15390_/Y VGND VGND VPWR VPWR _15398_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14342_ _15875_/A _14256_/B _14256_/Y VGND VGND VPWR VPWR _14342_/Y sky130_fd_sc_hd__o21ai_1
X_11554_ _11488_/Y _11553_/Y _11488_/Y _11553_/Y VGND VGND VPWR VPWR _11557_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14273_ _14273_/A VGND VGND VPWR VPWR _14273_/Y sky130_fd_sc_hd__inv_2
X_10505_ _13605_/A _10527_/B VGND VGND VPWR VPWR _10505_/Y sky130_fd_sc_hd__nor2_1
X_11485_ _09439_/X _11484_/X _09439_/X _11484_/X VGND VGND VPWR VPWR _11486_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16012_ _15955_/X _16011_/Y _15955_/X _16011_/Y VGND VGND VPWR VPWR _16038_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13224_ _13201_/X _13223_/Y _13201_/X _13223_/Y VGND VGND VPWR VPWR _13300_/B sky130_fd_sc_hd__a2bb2o_1
X_10436_ _09312_/A _09312_/B _09312_/Y VGND VGND VPWR VPWR _10438_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13155_ _13116_/X _13154_/Y _13116_/X _13154_/Y VGND VGND VPWR VPWR _13198_/B sky130_fd_sc_hd__a2bb2o_1
X_10367_ _10367_/A _11753_/A VGND VGND VPWR VPWR _10367_/Y sky130_fd_sc_hd__nor2_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12106_ _12106_/A _12157_/B VGND VGND VPWR VPWR _12106_/Y sky130_fd_sc_hd__nand2_1
X_13086_ _13016_/X _13085_/X _13016_/X _13085_/X VGND VGND VPWR VPWR _13107_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10325_/A _12702_/A VGND VGND VPWR VPWR _10298_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12037_ _11968_/A _11968_/B _11968_/Y VGND VGND VPWR VPWR _12037_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13988_ _13988_/A _13988_/B VGND VGND VPWR VPWR _13988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15727_ _14921_/X _15726_/X _14921_/X _15726_/X VGND VGND VPWR VPWR _15728_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12939_ _12888_/Y _12937_/X _12938_/Y VGND VGND VPWR VPWR _12939_/X sky130_fd_sc_hd__o21a_1
X_15658_ _15658_/A VGND VGND VPWR VPWR _15658_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14609_ _15347_/A _14661_/B VGND VGND VPWR VPWR _14609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15589_ _16046_/A VGND VGND VPWR VPWR _15683_/A sky130_fd_sc_hd__inv_2
XFILLER_103_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08963_ _08962_/X _10125_/A _08827_/Y VGND VGND VPWR VPWR _08963_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08894_ _08893_/X _08793_/B _08793_/Y VGND VGND VPWR VPWR _08894_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09515_ _09486_/A _09486_/B _09486_/Y _09514_/X VGND VGND VPWR VPWR _09515_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09446_ _09247_/A _09428_/A _09262_/A _09428_/Y _10929_/A VGND VGND VPWR VPWR _12065_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_25_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09377_ _09472_/B _09860_/A _09352_/A VGND VGND VPWR VPWR _09377_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08328_ _08328_/A VGND VGND VPWR VPWR _08328_/Y sky130_fd_sc_hd__inv_2
X_08259_ input31/X VGND VGND VPWR VPWR _08260_/B sky130_fd_sc_hd__inv_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11270_ _09431_/B _09376_/B _09376_/X VGND VGND VPWR VPWR _11271_/B sky130_fd_sc_hd__a21boi_1
XFILLER_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10221_ _10180_/A _10180_/B _10180_/Y VGND VGND VPWR VPWR _10222_/A sky130_fd_sc_hd__o21ai_1
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10152_ _10116_/A _10116_/B _10117_/A VGND VGND VPWR VPWR _10155_/A sky130_fd_sc_hd__a21bo_1
XFILLER_94_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14960_ _14957_/X _14959_/X _14957_/X _14959_/X VGND VGND VPWR VPWR _14971_/B sky130_fd_sc_hd__a2bb2o_1
X_10083_ _10083_/A _10083_/B VGND VGND VPWR VPWR _11142_/B sky130_fd_sc_hd__or2_1
XFILLER_102_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13911_ _13848_/X _13910_/Y _13848_/X _13910_/Y VGND VGND VPWR VPWR _13949_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14891_ _14819_/X _14890_/X _14819_/X _14890_/X VGND VGND VPWR VPWR _14912_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13842_ _13827_/Y _13840_/X _13841_/Y VGND VGND VPWR VPWR _13842_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13773_ _13803_/A _13771_/X _13772_/X VGND VGND VPWR VPWR _13773_/X sky130_fd_sc_hd__o21a_1
X_15512_ _15512_/A _15512_/B VGND VGND VPWR VPWR _15512_/X sky130_fd_sc_hd__and2_1
X_12724_ _13457_/A _13457_/B _12723_/Y VGND VGND VPWR VPWR _12724_/Y sky130_fd_sc_hd__o21ai_1
X_10985_ _10983_/A _10983_/B _10983_/Y _10984_/X VGND VGND VPWR VPWR _12174_/A sky130_fd_sc_hd__o211a_1
XFILLER_31_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15443_ _15443_/A _15443_/B VGND VGND VPWR VPWR _15443_/X sky130_fd_sc_hd__and2_1
X_12655_ _13978_/A VGND VGND VPWR VPWR _14948_/A sky130_fd_sc_hd__inv_2
XFILLER_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12586_ _12586_/A VGND VGND VPWR VPWR _12586_/Y sky130_fd_sc_hd__inv_2
X_15374_ _15410_/A _15410_/B VGND VGND VPWR VPWR _15450_/A sky130_fd_sc_hd__and2_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11606_ _10088_/X _11605_/X _10088_/X _11605_/X VGND VGND VPWR VPWR _11607_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14325_ _14264_/A _14324_/Y _14264_/A _14324_/Y VGND VGND VPWR VPWR _14387_/A sky130_fd_sc_hd__a2bb2o_1
X_11537_ _11536_/A _11536_/B _11536_/Y _10984_/X VGND VGND VPWR VPWR _12419_/A sky130_fd_sc_hd__o211a_2
X_14256_ _15875_/A _14256_/B VGND VGND VPWR VPWR _14256_/Y sky130_fd_sc_hd__nand2_1
X_11468_ _15440_/A _11355_/B _11355_/Y _11263_/X VGND VGND VPWR VPWR _11468_/X sky130_fd_sc_hd__a2bb2o_1
X_14187_ _14115_/X _14186_/Y _14115_/X _14186_/Y VGND VGND VPWR VPWR _14188_/B sky130_fd_sc_hd__a2bb2oi_1
X_13207_ _13144_/Y _13205_/X _13206_/Y VGND VGND VPWR VPWR _13207_/X sky130_fd_sc_hd__o21a_1
X_10419_ _10354_/X _10418_/Y _10354_/X _10418_/Y VGND VGND VPWR VPWR _10429_/B sky130_fd_sc_hd__a2bb2o_1
X_11399_ _11399_/A VGND VGND VPWR VPWR _11399_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13138_ _13126_/X _13137_/Y _13126_/X _13137_/Y VGND VGND VPWR VPWR _13139_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _13766_/A VGND VGND VPWR VPWR _15252_/A sky130_fd_sc_hd__buf_1
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09300_ _09300_/A VGND VGND VPWR VPWR _09300_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09231_ _09540_/A _09684_/A VGND VGND VPWR VPWR _09231_/Y sky130_fd_sc_hd__nor2_1
X_09162_ _08749_/Y _09161_/Y _08749_/Y _09161_/Y VGND VGND VPWR VPWR _10008_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09093_ _10017_/B _09072_/B _09073_/B VGND VGND VPWR VPWR _09705_/A sky130_fd_sc_hd__a21bo_1
XFILLER_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09995_ _09995_/A _09995_/B VGND VGND VPWR VPWR _11308_/B sky130_fd_sc_hd__or2_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08946_ _08946_/A VGND VGND VPWR VPWR _08946_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08877_ _08691_/X _08876_/Y _08691_/X _08876_/Y VGND VGND VPWR VPWR _08982_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10770_ _10904_/A _10767_/X _10769_/X VGND VGND VPWR VPWR _10770_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09429_ _09429_/A _09429_/B VGND VGND VPWR VPWR _09429_/X sky130_fd_sc_hd__or2_1
XFILLER_100_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12440_ _12439_/A _12439_/B _12439_/X VGND VGND VPWR VPWR _12441_/B sky130_fd_sc_hd__a21bo_1
XFILLER_126_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14110_ _14053_/X _14109_/X _14053_/X _14109_/X VGND VGND VPWR VPWR _14110_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12371_ _12371_/A _12371_/B VGND VGND VPWR VPWR _12371_/X sky130_fd_sc_hd__or2_1
X_15090_ _15081_/A _15081_/B _15081_/Y _15089_/X VGND VGND VPWR VPWR _15090_/X sky130_fd_sc_hd__a2bb2o_1
X_11322_ _10239_/B _10143_/B _10143_/Y VGND VGND VPWR VPWR _11323_/A sky130_fd_sc_hd__a21oi_1
X_11253_ _11250_/X _11251_/X _11419_/B VGND VGND VPWR VPWR _11253_/X sky130_fd_sc_hd__o21a_1
X_14041_ _13938_/X _14040_/X _13938_/X _14040_/X VGND VGND VPWR VPWR _14042_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10204_ _08664_/X _09404_/Y _08671_/A _09403_/X VGND VGND VPWR VPWR _10902_/B sky130_fd_sc_hd__o22a_2
XFILLER_121_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11184_ _14014_/A VGND VGND VPWR VPWR _14059_/A sky130_fd_sc_hd__buf_1
X_15992_ _15990_/X _15992_/B VGND VGND VPWR VPWR _15992_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10135_ _10134_/A _10134_/B _10134_/X VGND VGND VPWR VPWR _10194_/A sky130_fd_sc_hd__a21bo_1
XFILLER_125_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14943_ _15425_/A _14980_/B _14942_/Y VGND VGND VPWR VPWR _14943_/Y sky130_fd_sc_hd__o21ai_1
X_10066_ _10021_/X _10065_/Y _10021_/X _10065_/Y VGND VGND VPWR VPWR _10067_/B sky130_fd_sc_hd__a2bb2o_1
X_14874_ _14824_/X _14873_/X _14824_/X _14873_/X VGND VGND VPWR VPWR _14922_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13825_ _13825_/A _13758_/X VGND VGND VPWR VPWR _13825_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13756_ _13756_/A _13756_/B VGND VGND VPWR VPWR _13756_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10968_ _10968_/A VGND VGND VPWR VPWR _11607_/A sky130_fd_sc_hd__clkbuf_2
X_13687_ _13679_/Y _13685_/Y _13686_/Y VGND VGND VPWR VPWR _13687_/X sky130_fd_sc_hd__o21a_1
X_12707_ _12707_/A _12707_/B VGND VGND VPWR VPWR _12707_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12638_ _12638_/A _12638_/B VGND VGND VPWR VPWR _12638_/X sky130_fd_sc_hd__or2_1
X_10899_ _10899_/A _10772_/X VGND VGND VPWR VPWR _10899_/X sky130_fd_sc_hd__or2b_1
X_15426_ _15159_/Y _15425_/Y _15171_/Y VGND VGND VPWR VPWR _15426_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12569_ _12569_/A VGND VGND VPWR VPWR _12569_/Y sky130_fd_sc_hd__inv_2
X_15357_ _15293_/X _15357_/B VGND VGND VPWR VPWR _15357_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14308_ _14308_/A _14308_/B VGND VGND VPWR VPWR _15964_/A sky130_fd_sc_hd__or2_1
X_15288_ _15284_/Y _15287_/Y _15284_/Y _15287_/Y VGND VGND VPWR VPWR _15289_/B sky130_fd_sc_hd__o2bb2a_1
X_14239_ _14239_/A VGND VGND VPWR VPWR _14243_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08800_ _09213_/A VGND VGND VPWR VPWR _10014_/A sky130_fd_sc_hd__buf_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _10081_/A _09778_/Y _09779_/Y VGND VGND VPWR VPWR _09782_/B sky130_fd_sc_hd__o21ai_2
XFILLER_79_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08731_ _08714_/Y _08729_/Y _08730_/X VGND VGND VPWR VPWR _08731_/Y sky130_fd_sc_hd__o21ai_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08662_ _08662_/A _08662_/B VGND VGND VPWR VPWR _09677_/A sky130_fd_sc_hd__or2_1
XFILLER_93_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08593_ _08592_/Y _08423_/X _08592_/Y _08423_/X VGND VGND VPWR VPWR _08596_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09214_ _09856_/A VGND VGND VPWR VPWR _09728_/A sky130_fd_sc_hd__inv_2
XFILLER_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09145_ _09145_/A VGND VGND VPWR VPWR _09145_/Y sky130_fd_sc_hd__inv_2
X_09076_ _10013_/B _09076_/B VGND VGND VPWR VPWR _09077_/B sky130_fd_sc_hd__or2_1
XFILLER_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09978_ _09978_/A _09978_/B VGND VGND VPWR VPWR _09978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08929_ _08929_/A _08929_/B VGND VGND VPWR VPWR _10287_/A sky130_fd_sc_hd__or2_1
X_11940_ _13698_/A _11980_/B _11939_/Y VGND VGND VPWR VPWR _11940_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11871_ _11870_/A _11912_/B _11870_/Y VGND VGND VPWR VPWR _11871_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14590_ _14522_/X _14536_/A _14535_/X VGND VGND VPWR VPWR _14590_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13610_ _12917_/Y _12918_/X _12917_/A _12916_/Y VGND VGND VPWR VPWR _13611_/A sky130_fd_sc_hd__a22o_1
XFILLER_60_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10822_ _10822_/A VGND VGND VPWR VPWR _10822_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10753_ _13756_/A VGND VGND VPWR VPWR _11966_/A sky130_fd_sc_hd__inv_2
XFILLER_53_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13541_ _15051_/A _13500_/B _13500_/Y _13540_/X VGND VGND VPWR VPWR _13541_/X sky130_fd_sc_hd__a2bb2o_1
X_16260_ _16260_/A _16260_/B VGND VGND VPWR VPWR _16260_/Y sky130_fd_sc_hd__nand2_1
X_13472_ _14367_/A VGND VGND VPWR VPWR _14352_/A sky130_fd_sc_hd__clkbuf_2
X_15211_ _15211_/A _15211_/B VGND VGND VPWR VPWR _15211_/Y sky130_fd_sc_hd__nand2_1
X_10684_ _10684_/A VGND VGND VPWR VPWR _10684_/Y sky130_fd_sc_hd__inv_2
X_16191_ _15808_/X _16190_/X _15808_/X _16190_/X VGND VGND VPWR VPWR _16192_/B sky130_fd_sc_hd__a2bb2o_1
X_12423_ _12422_/A _12422_/B _12422_/Y VGND VGND VPWR VPWR _12435_/B sky130_fd_sc_hd__o21ai_2
X_12354_ _12311_/A _12311_/B _12311_/Y _12535_/A VGND VGND VPWR VPWR _12527_/A sky130_fd_sc_hd__a2bb2o_1
X_15142_ _15088_/X _15141_/Y _15088_/X _15141_/Y VGND VGND VPWR VPWR _15143_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15073_ _15073_/A _15034_/X VGND VGND VPWR VPWR _15073_/X sky130_fd_sc_hd__or2b_1
X_11305_ _11304_/A _11304_/B _11304_/X _11129_/X VGND VGND VPWR VPWR _11305_/X sky130_fd_sc_hd__o22a_1
X_14024_ _14027_/A VGND VGND VPWR VPWR _15458_/A sky130_fd_sc_hd__buf_1
X_12285_ _12260_/X _12284_/Y _12260_/X _12284_/Y VGND VGND VPWR VPWR _12364_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11236_ _11236_/A _11080_/X VGND VGND VPWR VPWR _11236_/X sky130_fd_sc_hd__or2b_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11167_ _12256_/A _11290_/B VGND VGND VPWR VPWR _11167_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10118_ _10118_/A _10118_/B VGND VGND VPWR VPWR _10119_/A sky130_fd_sc_hd__or2_1
X_15975_ _14162_/X _15853_/A _14162_/X _15853_/A VGND VGND VPWR VPWR _15984_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11098_ _11097_/A _11097_/B _11097_/Y _09392_/X VGND VGND VPWR VPWR _11304_/A sky130_fd_sc_hd__o211a_1
XFILLER_36_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14926_ _15550_/A _14926_/B VGND VGND VPWR VPWR _14926_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10049_ _10049_/A _10079_/B VGND VGND VPWR VPWR _10049_/X sky130_fd_sc_hd__and2_1
XFILLER_90_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14857_ _14858_/A _14858_/B VGND VGND VPWR VPWR _14859_/A sky130_fd_sc_hd__and2_1
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14788_ _14788_/A _14734_/X VGND VGND VPWR VPWR _14788_/X sky130_fd_sc_hd__or2b_1
X_13808_ _14610_/A _13853_/B VGND VGND VPWR VPWR _13808_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13739_ _13691_/X _13738_/X _13691_/X _13738_/X VGND VGND VPWR VPWR _13762_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16458_ _16357_/A _16458_/D VGND VGND VPWR VPWR _16458_/Q sky130_fd_sc_hd__dfxtp_1
X_16389_ _16385_/X _16388_/Y _16385_/X _16388_/Y VGND VGND VPWR VPWR _16389_/X sky130_fd_sc_hd__a2bb2o_1
X_15409_ _15453_/A _15407_/X _15408_/X VGND VGND VPWR VPWR _15409_/X sky130_fd_sc_hd__o21a_1
XFILLER_117_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09901_ _09898_/X _09901_/B VGND VGND VPWR VPWR _09903_/B sky130_fd_sc_hd__nand2b_1
XFILLER_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09832_ _09832_/A _09832_/B VGND VGND VPWR VPWR _09833_/A sky130_fd_sc_hd__nand2_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _09763_/A VGND VGND VPWR VPWR _09779_/A sky130_fd_sc_hd__inv_2
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08714_ _08714_/A _08714_/B VGND VGND VPWR VPWR _08714_/Y sky130_fd_sc_hd__nor2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _08605_/X _09696_/B _08605_/X _09696_/B VGND VGND VPWR VPWR _09695_/B sky130_fd_sc_hd__a2bb2o_1
Xrebuffer10 rebuffer11/X VGND VGND VPWR VPWR rebuffer9/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer21 _10194_/B VGND VGND VPWR VPWR rebuffer21/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer54 _10206_/A VGND VGND VPWR VPWR _12657_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_08645_ _08645_/A VGND VGND VPWR VPWR _08645_/X sky130_fd_sc_hd__buf_1
Xrebuffer43 _09749_/X VGND VGND VPWR VPWR _10001_/B1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer32 _10173_/A VGND VGND VPWR VPWR _10248_/A sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _08589_/A _08576_/B VGND VGND VPWR VPWR _09454_/B sky130_fd_sc_hd__or2_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09128_ _09424_/A _09131_/B VGND VGND VPWR VPWR _09128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09059_ _08806_/Y _09047_/A _08806_/A _09047_/Y VGND VGND VPWR VPWR _10015_/B sky130_fd_sc_hd__o22a_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12070_ _12070_/A _12070_/B VGND VGND VPWR VPWR _12070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11021_ _10920_/X _11020_/X _10920_/X _11020_/X VGND VGND VPWR VPWR _11090_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15760_ _14910_/A _14910_/B _14910_/Y VGND VGND VPWR VPWR _15760_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12972_ _13700_/A VGND VGND VPWR VPWR _14523_/A sky130_fd_sc_hd__inv_2
XFILLER_58_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15691_ _15549_/X _15690_/X _15549_/X _15690_/X VGND VGND VPWR VPWR _15692_/B sky130_fd_sc_hd__a2bb2o_1
X_14711_ _15333_/A _14647_/B _14647_/Y VGND VGND VPWR VPWR _14711_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11923_ _11923_/A _11923_/B VGND VGND VPWR VPWR _11923_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14642_ _13096_/X _14641_/Y _13096_/X _14641_/Y VGND VGND VPWR VPWR _14643_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11854_ _11916_/A VGND VGND VPWR VPWR _12774_/A sky130_fd_sc_hd__buf_1
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10805_ _13512_/A _10804_/B _10804_/X _10668_/X VGND VGND VPWR VPWR _10805_/X sky130_fd_sc_hd__o22a_1
X_14573_ _15272_/A _14573_/B VGND VGND VPWR VPWR _14573_/Y sky130_fd_sc_hd__nand2_1
X_11785_ _11790_/A VGND VGND VPWR VPWR _14428_/A sky130_fd_sc_hd__buf_1
XFILLER_41_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16312_ _16457_/X VGND VGND VPWR VPWR _16312_/Y sky130_fd_sc_hd__inv_4
X_13524_ _13524_/A _13524_/B VGND VGND VPWR VPWR _13524_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10736_ _10736_/A VGND VGND VPWR VPWR _10736_/Y sky130_fd_sc_hd__inv_2
X_16243_ _16243_/A _16384_/B VGND VGND VPWR VPWR _16244_/A sky130_fd_sc_hd__or2_1
X_13455_ _13453_/X _13454_/Y _13453_/X _13454_/Y VGND VGND VPWR VPWR _13455_/X sky130_fd_sc_hd__a2bb2o_1
X_10667_ _11853_/A _10667_/B VGND VGND VPWR VPWR _10667_/X sky130_fd_sc_hd__and2_1
XFILLER_127_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16174_ _16112_/A _15813_/B _15813_/Y VGND VGND VPWR VPWR _16174_/X sky130_fd_sc_hd__o21a_1
X_12406_ _12359_/X _12405_/Y _12359_/X _12405_/Y VGND VGND VPWR VPWR _12407_/B sky130_fd_sc_hd__a2bb2o_1
X_13386_ _14125_/A _13441_/B VGND VGND VPWR VPWR _13386_/Y sky130_fd_sc_hd__nor2_1
X_15125_ _15125_/A _15125_/B VGND VGND VPWR VPWR _15125_/Y sky130_fd_sc_hd__nand2_1
X_10598_ _10598_/A VGND VGND VPWR VPWR _10598_/Y sky130_fd_sc_hd__inv_2
X_12337_ _12333_/Y _12581_/A _12336_/Y VGND VGND VPWR VPWR _12341_/B sky130_fd_sc_hd__o21ai_1
XFILLER_126_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15056_ _15045_/X _15055_/X _15045_/X _15055_/X VGND VGND VPWR VPWR _15057_/B sky130_fd_sc_hd__a2bb2o_1
X_12268_ _12268_/A _12268_/B VGND VGND VPWR VPWR _12268_/X sky130_fd_sc_hd__or2_1
X_11219_ _12220_/A _11219_/B VGND VGND VPWR VPWR _11219_/Y sky130_fd_sc_hd__nand2_1
X_14007_ _13958_/X _14006_/Y _13958_/X _14006_/Y VGND VGND VPWR VPWR _14063_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12199_ _13202_/A _12251_/B _12198_/Y VGND VGND VPWR VPWR _12199_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15958_ _15958_/A _15958_/B VGND VGND VPWR VPWR _16008_/B sky130_fd_sc_hd__or2_1
XFILLER_76_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14909_ _14898_/Y _14907_/X _14908_/Y VGND VGND VPWR VPWR _14909_/X sky130_fd_sc_hd__o21a_1
X_15889_ _15880_/Y _15887_/X _15888_/Y VGND VGND VPWR VPWR _15889_/X sky130_fd_sc_hd__o21a_1
X_08430_ _08429_/A _08333_/Y _08429_/Y _08333_/A _08441_/A VGND VGND VPWR VPWR _09209_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08361_ _08361_/A VGND VGND VPWR VPWR _08361_/Y sky130_fd_sc_hd__inv_2
X_08292_ _08321_/A input19/X _08322_/A _08324_/A VGND VGND VPWR VPWR _08319_/A sky130_fd_sc_hd__o22a_1
XFILLER_32_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09815_ _09810_/X _08830_/A _09810_/X _08830_/A VGND VGND VPWR VPWR _09819_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09746_ _09347_/B _09743_/X _08512_/X VGND VGND VPWR VPWR _09791_/B sky130_fd_sc_hd__o21a_1
XFILLER_27_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09677_/A _09677_/B VGND VGND VPWR VPWR _09681_/B sky130_fd_sc_hd__and2_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08628_ _08634_/A VGND VGND VPWR VPWR _09458_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08559_ _08558_/A _08439_/Y _08558_/Y _08439_/A VGND VGND VPWR VPWR _10117_/B sky130_fd_sc_hd__o22a_1
X_11570_ _08986_/A _08986_/B _08986_/Y VGND VGND VPWR VPWR _11570_/X sky130_fd_sc_hd__o21a_1
X_10521_ _10521_/A _10625_/C VGND VGND VPWR VPWR _10522_/A sky130_fd_sc_hd__or2_1
XFILLER_10_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13240_ _14734_/A _13291_/B VGND VGND VPWR VPWR _13240_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10452_ _11808_/A _10452_/B VGND VGND VPWR VPWR _10452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13171_ _13188_/A _13188_/B VGND VGND VPWR VPWR _13171_/Y sky130_fd_sc_hd__nor2_1
X_10383_ _10252_/A _10252_/B _10252_/Y VGND VGND VPWR VPWR _10384_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12122_ _13190_/A _12057_/B _12057_/Y VGND VGND VPWR VPWR _12122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12053_ _12053_/A _12053_/B VGND VGND VPWR VPWR _12053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11004_ _11004_/A VGND VGND VPWR VPWR _14409_/A sky130_fd_sc_hd__buf_1
X_15812_ _15743_/Y _15810_/X _15811_/Y VGND VGND VPWR VPWR _15812_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15743_ _16110_/A _15811_/B VGND VGND VPWR VPWR _15743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12955_ _12955_/A VGND VGND VPWR VPWR _13878_/A sky130_fd_sc_hd__inv_2
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11906_ _11906_/A VGND VGND VPWR VPWR _11906_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15674_ _15630_/Y _15672_/X _15673_/Y VGND VGND VPWR VPWR _15674_/X sky130_fd_sc_hd__o21a_1
XFILLER_73_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12886_ _12851_/A _12851_/B _12851_/Y VGND VGND VPWR VPWR _12886_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _15339_/A _14653_/B VGND VGND VPWR VPWR _14625_/Y sky130_fd_sc_hd__nor2_1
X_11837_ _13609_/A _11836_/B _10626_/A _11836_/Y VGND VGND VPWR VPWR _11837_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14556_/A _14513_/X VGND VGND VPWR VPWR _14556_/X sky130_fd_sc_hd__or2b_1
X_11768_ _11766_/X _11768_/B VGND VGND VPWR VPWR _11768_/Y sky130_fd_sc_hd__nand2b_1
X_13507_ _13509_/A VGND VGND VPWR VPWR _15042_/A sky130_fd_sc_hd__buf_1
XFILLER_41_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10719_ _10933_/A _10719_/B VGND VGND VPWR VPWR _13073_/A sky130_fd_sc_hd__or2_2
X_14487_ _15199_/A _14517_/B VGND VGND VPWR VPWR _14548_/A sky130_fd_sc_hd__and2_1
X_11699_ _11695_/Y _11698_/X _11695_/Y _11698_/X VGND VGND VPWR VPWR _11699_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16226_ _16094_/A _15795_/B _15795_/Y VGND VGND VPWR VPWR _16228_/A sky130_fd_sc_hd__o21ai_1
X_13438_ _13392_/Y _13436_/X _13437_/Y VGND VGND VPWR VPWR _13438_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer1 rebuffer3/X VGND VGND VPWR VPWR _11609_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_16157_ _16388_/A _16157_/B VGND VGND VPWR VPWR _16268_/A sky130_fd_sc_hd__or2_1
X_13369_ _13381_/A _13367_/X _13368_/X VGND VGND VPWR VPWR _13369_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16088_ _16029_/X _16087_/Y _16029_/X _16087_/Y VGND VGND VPWR VPWR _16223_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15108_ _15107_/A _15107_/B _15107_/Y VGND VGND VPWR VPWR _15108_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15039_ _15067_/A _15037_/X _15038_/X VGND VGND VPWR VPWR _15039_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09600_ _09983_/A VGND VGND VPWR VPWR _09984_/A sky130_fd_sc_hd__buf_1
X_09531_ _09531_/A _09531_/B VGND VGND VPWR VPWR _09532_/A sky130_fd_sc_hd__or2_1
XFILLER_83_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09462_ _10018_/A _09462_/B VGND VGND VPWR VPWR _09462_/X sky130_fd_sc_hd__or2_1
X_09393_ _09329_/A _09329_/B _09329_/Y _09392_/X VGND VGND VPWR VPWR _11128_/A sky130_fd_sc_hd__o211a_1
XFILLER_12_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08413_ _09225_/B _08408_/Y _09251_/A VGND VGND VPWR VPWR _08413_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08344_ _08344_/A VGND VGND VPWR VPWR _08344_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08275_ _08275_/A input10/X VGND VGND VPWR VPWR _08387_/A sky130_fd_sc_hd__nor2_1
XFILLER_118_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09729_ _08580_/X _09731_/B _08580_/X _09731_/B VGND VGND VPWR VPWR _09730_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ _12693_/A _12693_/B _12693_/Y VGND VGND VPWR VPWR _12740_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A VGND VGND VPWR VPWR _12671_/Y sky130_fd_sc_hd__inv_2
X_15390_ _15331_/A _15331_/B _15331_/Y VGND VGND VPWR VPWR _15390_/Y sky130_fd_sc_hd__o21ai_1
X_14410_ _15246_/A VGND VGND VPWR VPWR _14587_/A sky130_fd_sc_hd__buf_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _12419_/A VGND VGND VPWR VPWR _12382_/A sky130_fd_sc_hd__inv_2
X_14341_ _14383_/A _15954_/A VGND VGND VPWR VPWR _14341_/X sky130_fd_sc_hd__and2_1
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11553_ _13882_/A _11652_/B _11552_/Y VGND VGND VPWR VPWR _11553_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14272_ _14191_/Y _14270_/Y _14271_/Y VGND VGND VPWR VPWR _14273_/A sky130_fd_sc_hd__o21ai_2
XFILLER_109_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10504_ _10432_/X _10503_/X _10432_/X _10503_/X VGND VGND VPWR VPWR _10527_/B sky130_fd_sc_hd__a2bb2o_1
X_11484_ _09788_/A _09367_/A _09430_/X VGND VGND VPWR VPWR _11484_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16011_ _15933_/X _16011_/B VGND VGND VPWR VPWR _16011_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13223_ _13202_/A _13202_/B _13202_/Y VGND VGND VPWR VPWR _13223_/Y sky130_fd_sc_hd__o21ai_1
X_10435_ _13559_/A _10392_/B _10392_/X _10434_/X VGND VGND VPWR VPWR _10435_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13154_ _15246_/A _13117_/B _13117_/Y VGND VGND VPWR VPWR _13154_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12105_ _12069_/X _12104_/Y _12069_/X _12104_/Y VGND VGND VPWR VPWR _12157_/B sky130_fd_sc_hd__a2bb2o_1
X_10366_ _11760_/A VGND VGND VPWR VPWR _11753_/A sky130_fd_sc_hd__clkinvlp_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13085_/A _13017_/X VGND VGND VPWR VPWR _13085_/X sky130_fd_sc_hd__or2b_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _10325_/B VGND VGND VPWR VPWR _12702_/A sky130_fd_sc_hd__inv_2
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12036_ _13188_/A _12055_/B VGND VGND VPWR VPWR _12036_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13987_ _13985_/Y _13986_/X _13985_/Y _13986_/X VGND VGND VPWR VPWR _13988_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15726_ _15546_/A _14922_/B _14922_/Y VGND VGND VPWR VPWR _15726_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12938_ _12938_/A _12938_/B VGND VGND VPWR VPWR _12938_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15657_ _15509_/A _15509_/B _15510_/A VGND VGND VPWR VPWR _15658_/A sky130_fd_sc_hd__o21ai_1
XFILLER_61_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14608_ _14588_/X _14607_/Y _14588_/X _14607_/Y VGND VGND VPWR VPWR _14661_/B sky130_fd_sc_hd__a2bb2o_1
X_12869_ _12946_/A VGND VGND VPWR VPWR _14757_/A sky130_fd_sc_hd__buf_1
XFILLER_61_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15588_ _15700_/A _15588_/B VGND VGND VPWR VPWR _16046_/A sky130_fd_sc_hd__or2_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14539_ _15249_/A VGND VGND VPWR VPWR _14585_/A sky130_fd_sc_hd__buf_1
XFILLER_134_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16209_ _16207_/A _16208_/A _16207_/Y _16208_/Y _15832_/A VGND VGND VPWR VPWR _16255_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08962_ _10017_/A VGND VGND VPWR VPWR _08962_/X sky130_fd_sc_hd__buf_1
XFILLER_69_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08893_ _10013_/A VGND VGND VPWR VPWR _08893_/X sky130_fd_sc_hd__buf_1
XFILLER_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09514_ _09488_/A _09488_/B _09488_/Y _09513_/X VGND VGND VPWR VPWR _09514_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09445_ _09445_/A VGND VGND VPWR VPWR _10929_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09376_ _09431_/B _09376_/B VGND VGND VPWR VPWR _09376_/X sky130_fd_sc_hd__or2_1
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08327_ _08327_/A _08327_/B VGND VGND VPWR VPWR _08328_/A sky130_fd_sc_hd__or2_1
X_08258_ input15/X VGND VGND VPWR VPWR _08336_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10220_ _11748_/A VGND VGND VPWR VPWR _10224_/A sky130_fd_sc_hd__inv_2
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10151_ _10151_/A _10151_/B VGND VGND VPWR VPWR _10151_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10082_ _10046_/X _10080_/X _10969_/B VGND VGND VPWR VPWR _10082_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13910_ _14618_/A _13849_/B _13849_/Y VGND VGND VPWR VPWR _13910_/Y sky130_fd_sc_hd__o21ai_1
X_14890_ _14802_/A _14802_/B _14802_/A _14802_/B VGND VGND VPWR VPWR _14890_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13841_ _14634_/A _13841_/B VGND VGND VPWR VPWR _13841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13772_ _13772_/A _13772_/B VGND VGND VPWR VPWR _13772_/X sky130_fd_sc_hd__or2_1
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10984_ _10984_/A VGND VGND VPWR VPWR _10984_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15511_ _15509_/A _15509_/B _12610_/A _15510_/Y VGND VGND VPWR VPWR _15512_/B sky130_fd_sc_hd__o22a_1
X_12723_ _13457_/A _13457_/B VGND VGND VPWR VPWR _12723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15442_ _15415_/X _15441_/X _15415_/X _15441_/X VGND VGND VPWR VPWR _15443_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12654_ _13984_/A VGND VGND VPWR VPWR _14976_/A sky130_fd_sc_hd__buf_1
XFILLER_128_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12585_ _12622_/A _12622_/B VGND VGND VPWR VPWR _14219_/A sky130_fd_sc_hd__and2_1
X_15373_ _15342_/X _15372_/X _15342_/X _15372_/X VGND VGND VPWR VPWR _15410_/B sky130_fd_sc_hd__a2bb2o_1
X_11605_ _11605_/A1 _10034_/B _10034_/Y VGND VGND VPWR VPWR _11605_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14324_ _15866_/A _14265_/B _14265_/Y VGND VGND VPWR VPWR _14324_/Y sky130_fd_sc_hd__o21ai_1
X_11536_ _11536_/A _11536_/B VGND VGND VPWR VPWR _11536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14255_ _14255_/A VGND VGND VPWR VPWR _14255_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11467_ _14063_/A VGND VGND VPWR VPWR _15440_/A sky130_fd_sc_hd__buf_1
X_13206_ _13206_/A _13206_/B VGND VGND VPWR VPWR _13206_/Y sky130_fd_sc_hd__nand2_1
X_14186_ _13439_/A _14120_/A _14118_/Y VGND VGND VPWR VPWR _14186_/Y sky130_fd_sc_hd__a21oi_1
X_10418_ _12832_/A _10355_/B _10356_/A VGND VGND VPWR VPWR _10418_/Y sky130_fd_sc_hd__o21ai_1
X_11398_ _11395_/Y _11397_/Y _11395_/A _11397_/A _12606_/B VGND VGND VPWR VPWR _13395_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13137_ _14976_/A _13127_/B _13127_/Y VGND VGND VPWR VPWR _13137_/Y sky130_fd_sc_hd__o21ai_1
X_10349_ _10349_/A VGND VGND VPWR VPWR _10350_/B sky130_fd_sc_hd__inv_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13068_ _13068_/A VGND VGND VPWR VPWR _13766_/A sky130_fd_sc_hd__inv_2
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12019_ _11977_/X _12018_/Y _11977_/X _12018_/Y VGND VGND VPWR VPWR _12063_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15709_ _15728_/A _15709_/B VGND VGND VPWR VPWR _16123_/A sky130_fd_sc_hd__or2_1
XFILLER_81_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09230_ _09230_/A _09800_/A VGND VGND VPWR VPWR _09230_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09161_ _08708_/Y _09160_/Y _08746_/X VGND VGND VPWR VPWR _09161_/Y sky130_fd_sc_hd__o21ai_1
X_09092_ _09703_/A VGND VGND VPWR VPWR _09418_/A sky130_fd_sc_hd__buf_1
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09994_ _09966_/Y _09992_/Y _09993_/Y VGND VGND VPWR VPWR _11309_/A sky130_fd_sc_hd__o21ai_1
XFILLER_88_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08945_ _08844_/A _08842_/Y _08944_/X VGND VGND VPWR VPWR _08946_/A sky130_fd_sc_hd__o21ai_1
XFILLER_57_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08876_ _08876_/A _08876_/B VGND VGND VPWR VPWR _08876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09428_ _09428_/A VGND VGND VPWR VPWR _09428_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09359_ _09344_/X _09358_/X _09344_/X _09358_/X VGND VGND VPWR VPWR _09359_/X sky130_fd_sc_hd__a2bb2o_1
X_12370_ _11275_/A _12369_/B _12369_/X _12262_/X VGND VGND VPWR VPWR _12370_/X sky130_fd_sc_hd__o22a_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11321_ _11321_/A VGND VGND VPWR VPWR _11521_/A sky130_fd_sc_hd__inv_2
XFILLER_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11252_ _14047_/A _11252_/B VGND VGND VPWR VPWR _11419_/B sky130_fd_sc_hd__or2_1
X_14040_ _14040_/A _13939_/X VGND VGND VPWR VPWR _14040_/X sky130_fd_sc_hd__or2b_1
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11183_ _13366_/A VGND VGND VPWR VPWR _14014_/A sky130_fd_sc_hd__inv_2
XFILLER_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10203_ _10215_/A _11245_/A VGND VGND VPWR VPWR _10282_/A sky130_fd_sc_hd__or2_2
XFILLER_69_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10134_ _10134_/A _10134_/B VGND VGND VPWR VPWR _10134_/X sky130_fd_sc_hd__or2_1
X_15991_ _15991_/A _15991_/B VGND VGND VPWR VPWR _15992_/B sky130_fd_sc_hd__or2_1
XFILLER_95_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14942_ _15171_/A _14980_/B VGND VGND VPWR VPWR _14942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10065_ _10065_/A _10065_/B VGND VGND VPWR VPWR _10065_/Y sky130_fd_sc_hd__nor2_1
X_14873_ _14782_/A _14782_/B _14782_/A _14782_/B VGND VGND VPWR VPWR _14873_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13824_ _13824_/A VGND VGND VPWR VPWR _14634_/A sky130_fd_sc_hd__inv_2
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13755_ _13752_/A _13752_/B _13752_/Y _13754_/Y VGND VGND VPWR VPWR _13755_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10967_ _10966_/Y _10815_/X _10824_/Y VGND VGND VPWR VPWR _10967_/X sky130_fd_sc_hd__o21a_1
X_16474_ _16474_/D _16454_/Y VGND VGND VPWR VPWR _16474_/Q sky130_fd_sc_hd__dlxtn_1
X_10898_ _13828_/A VGND VGND VPWR VPWR _13184_/A sky130_fd_sc_hd__buf_1
X_13686_ _14500_/A _13686_/B VGND VGND VPWR VPWR _13686_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12706_ _12705_/Y _12657_/Y _12705_/Y _12657_/Y VGND VGND VPWR VPWR _12707_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12637_ _14177_/A _12635_/X _12636_/X VGND VGND VPWR VPWR _12637_/X sky130_fd_sc_hd__o21a_1
X_15425_ _15425_/A _15425_/B VGND VGND VPWR VPWR _15425_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12568_ _14912_/A _11443_/B _11443_/Y VGND VGND VPWR VPWR _12569_/A sky130_fd_sc_hd__o21ai_1
X_15356_ _15422_/A _15422_/B VGND VGND VPWR VPWR _15356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14307_ _13440_/X _14306_/X _13440_/X _14306_/X VGND VGND VPWR VPWR _14308_/B sky130_fd_sc_hd__a2bb2oi_1
X_12499_ _12475_/X _12498_/X _12475_/X _12498_/X VGND VGND VPWR VPWR _12649_/A sky130_fd_sc_hd__a2bb2o_4
X_15287_ _15287_/A _15287_/B VGND VGND VPWR VPWR _15287_/Y sky130_fd_sc_hd__nor2_1
X_11519_ _11519_/A _12275_/A VGND VGND VPWR VPWR _11519_/Y sky130_fd_sc_hd__nor2_1
X_14238_ _14238_/A VGND VGND VPWR VPWR _14238_/Y sky130_fd_sc_hd__clkinvlp_2
X_14169_ _14281_/A _14169_/B VGND VGND VPWR VPWR _15910_/A sky130_fd_sc_hd__or2_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08730_ _09213_/A _09454_/B VGND VGND VPWR VPWR _08730_/X sky130_fd_sc_hd__or2_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08661_ _08919_/A VGND VGND VPWR VPWR _09234_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08592_ _08592_/A VGND VGND VPWR VPWR _08592_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09213_ _09213_/A _09213_/B VGND VGND VPWR VPWR _09856_/A sky130_fd_sc_hd__or2_1
XFILLER_22_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09144_ _09432_/A _09175_/B _09143_/Y VGND VGND VPWR VPWR _09145_/A sky130_fd_sc_hd__o21ai_1
XFILLER_108_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09075_ _10014_/B _09075_/B VGND VGND VPWR VPWR _09076_/B sky130_fd_sc_hd__or2_1
XFILLER_122_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09977_ _09977_/A _09978_/B VGND VGND VPWR VPWR _09977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08928_ _08928_/A VGND VGND VPWR VPWR _08929_/B sky130_fd_sc_hd__inv_2
XFILLER_57_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08859_ _09500_/A _08834_/A _08836_/Y _08955_/A VGND VGND VPWR VPWR _08859_/X sky130_fd_sc_hd__o22a_1
XFILLER_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11870_ _11870_/A _11912_/B VGND VGND VPWR VPWR _11870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10821_ _10821_/A VGND VGND VPWR VPWR _10821_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13540_ _15046_/A _13503_/B _13503_/Y _13539_/X VGND VGND VPWR VPWR _13540_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10752_ _09635_/A _10751_/A _09635_/Y _10751_/Y _09672_/A VGND VGND VPWR VPWR _13756_/A
+ sky130_fd_sc_hd__a221o_2
X_13471_ _13456_/X _13470_/X _13456_/X _13470_/X VGND VGND VPWR VPWR _14367_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15210_ _15147_/X _15209_/Y _15147_/X _15209_/Y VGND VGND VPWR VPWR _15211_/B sky130_fd_sc_hd__a2bb2o_1
X_12422_ _12422_/A _12422_/B VGND VGND VPWR VPWR _12422_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10683_ _10243_/B _10159_/B _10159_/Y VGND VGND VPWR VPWR _10684_/A sky130_fd_sc_hd__a21oi_1
X_16190_ _16108_/A _15809_/B _15809_/Y VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__o21a_1
X_12353_ _12314_/A _12314_/B _12314_/Y _12543_/A VGND VGND VPWR VPWR _12535_/A sky130_fd_sc_hd__a2bb2o_1
X_15141_ _15084_/A _15084_/B _15084_/Y VGND VGND VPWR VPWR _15141_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15072_ _15072_/A _15072_/B VGND VGND VPWR VPWR _15072_/Y sky130_fd_sc_hd__nand2_1
X_12284_ _13788_/A _12367_/B _12283_/Y VGND VGND VPWR VPWR _12284_/Y sky130_fd_sc_hd__o21ai_1
X_11304_ _11304_/A _11304_/B VGND VGND VPWR VPWR _11304_/X sky130_fd_sc_hd__and2_1
XFILLER_5_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11235_ _14038_/A VGND VGND VPWR VPWR _13344_/A sky130_fd_sc_hd__buf_1
X_14023_ _14023_/A _14023_/B VGND VGND VPWR VPWR _14023_/X sky130_fd_sc_hd__and2_1
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11166_ _11123_/X _11165_/Y _11123_/X _11165_/Y VGND VGND VPWR VPWR _11290_/B sky130_fd_sc_hd__a2bb2o_1
X_15974_ _15974_/A VGND VGND VPWR VPWR _15984_/A sky130_fd_sc_hd__inv_2
XFILLER_95_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11097_ _11097_/A _11097_/B VGND VGND VPWR VPWR _11097_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10117_ _10117_/A _10117_/B VGND VGND VPWR VPWR _10118_/A sky130_fd_sc_hd__or2_1
X_14925_ _14871_/Y _14923_/X _14924_/Y VGND VGND VPWR VPWR _14925_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10048_ _10025_/X _10047_/Y _10025_/X _10047_/Y VGND VGND VPWR VPWR _10079_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14856_ _14831_/X _14855_/Y _14831_/X _14855_/Y VGND VGND VPWR VPWR _14858_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08231__1 _08229_/A VGND VGND VPWR VPWR _16358_/A sky130_fd_sc_hd__inv_2
X_14787_ _15452_/A VGND VGND VPWR VPWR _14790_/A sky130_fd_sc_hd__buf_1
XFILLER_90_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13807_ _13769_/X _13806_/X _13769_/X _13806_/X VGND VGND VPWR VPWR _13853_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13738_ _13738_/A _13692_/X VGND VGND VPWR VPWR _13738_/X sky130_fd_sc_hd__or2b_1
X_11999_ _11999_/A _11999_/B VGND VGND VPWR VPWR _12000_/B sky130_fd_sc_hd__or2_1
XFILLER_31_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16457_ _16395_/A _16248_/B _16457_/S VGND VGND VPWR VPWR _16457_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13669_ _13692_/A _13692_/B VGND VGND VPWR VPWR _13738_/A sky130_fd_sc_hd__and2_1
XFILLER_129_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16388_ _16388_/A _16388_/B VGND VGND VPWR VPWR _16388_/Y sky130_fd_sc_hd__nor2_1
X_15408_ _15408_/A _15408_/B VGND VGND VPWR VPWR _15408_/X sky130_fd_sc_hd__or2_1
XFILLER_117_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15339_ _15339_/A _15339_/B VGND VGND VPWR VPWR _15339_/X sky130_fd_sc_hd__or2_1
X_09900_ _09898_/A _09898_/B _09899_/Y VGND VGND VPWR VPWR _09901_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _09829_/A _09829_/B _09830_/Y _08931_/Y VGND VGND VPWR VPWR _09832_/B sky130_fd_sc_hd__o22a_1
XFILLER_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _10046_/A VGND VGND VPWR VPWR _10081_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08713_/A _08713_/B VGND VGND VPWR VPWR _08713_/X sky130_fd_sc_hd__or2_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09693_ _09693_/A _09693_/B VGND VGND VPWR VPWR _09696_/B sky130_fd_sc_hd__or2_1
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer11 rebuffer12/X VGND VGND VPWR VPWR rebuffer11/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer55 _10206_/A VGND VGND VPWR VPWR _10283_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer33 _10248_/A VGND VGND VPWR VPWR _10314_/A1 sky130_fd_sc_hd__dlygate4sd1_1
X_08644_ _09458_/A _09228_/B _09228_/A _08386_/Y VGND VGND VPWR VPWR _08645_/A sky130_fd_sc_hd__o22a_1
XFILLER_27_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer44 _10001_/B1 VGND VGND VPWR VPWR _09790_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer22 _10191_/X VGND VGND VPWR VPWR rebuffer22/X sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08575_ _08574_/A _08338_/Y _08574_/Y _08338_/A VGND VGND VPWR VPWR _08576_/B sky130_fd_sc_hd__o22a_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09127_ _09088_/Y _09125_/Y _09126_/Y VGND VGND VPWR VPWR _09131_/B sky130_fd_sc_hd__o21ai_1
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09058_ _08798_/X _09048_/Y _08798_/X _09048_/Y VGND VGND VPWR VPWR _10014_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11020_ _11020_/A _10922_/X VGND VGND VPWR VPWR _11020_/X sky130_fd_sc_hd__or2b_1
XFILLER_2_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12971_ _14591_/A _13029_/B VGND VGND VPWR VPWR _13055_/A sky130_fd_sc_hd__and2_1
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15690_ _15494_/X _15690_/B VGND VGND VPWR VPWR _15690_/X sky130_fd_sc_hd__and2b_1
X_14710_ _14726_/A _14726_/B VGND VGND VPWR VPWR _14804_/A sky130_fd_sc_hd__and2_1
XFILLER_85_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11922_ _11921_/A _11921_/B _11921_/X _11862_/B VGND VGND VPWR VPWR _11992_/B sky130_fd_sc_hd__a22o_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14641_ _15270_/A _14571_/B _14571_/Y VGND VGND VPWR VPWR _14641_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11853_ _11853_/A VGND VGND VPWR VPWR _11916_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_45_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10804_ _11919_/A _10804_/B VGND VGND VPWR VPWR _10804_/X sky130_fd_sc_hd__and2_1
XFILLER_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16311_ _16318_/A _16318_/B VGND VGND VPWR VPWR _16311_/Y sky130_fd_sc_hd__nor2_1
X_14572_ _13096_/X _14570_/Y _14571_/Y VGND VGND VPWR VPWR _14572_/X sky130_fd_sc_hd__o21a_1
X_11784_ _12826_/A VGND VGND VPWR VPWR _11790_/A sky130_fd_sc_hd__inv_2
X_13523_ _10317_/X _13482_/X _10317_/X _13482_/X VGND VGND VPWR VPWR _13524_/B sky130_fd_sc_hd__o2bb2a_1
X_10735_ _10735_/A VGND VGND VPWR VPWR _10735_/Y sky130_fd_sc_hd__inv_2
X_16242_ _15784_/A _15784_/B _16241_/Y VGND VGND VPWR VPWR _16384_/B sky130_fd_sc_hd__a21oi_1
X_13454_ _14067_/A _13309_/B _13309_/Y _13372_/X VGND VGND VPWR VPWR _13454_/Y sky130_fd_sc_hd__o2bb2ai_1
X_10666_ _11016_/A VGND VGND VPWR VPWR _10666_/X sky130_fd_sc_hd__buf_1
X_16173_ _16189_/A _16173_/B VGND VGND VPWR VPWR _16264_/A sky130_fd_sc_hd__or2_1
X_13385_ _13365_/X _13384_/X _13365_/X _13384_/X VGND VGND VPWR VPWR _13441_/B sky130_fd_sc_hd__a2bb2o_1
X_12405_ _12403_/X _12405_/B VGND VGND VPWR VPWR _12405_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_127_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15124_ _15094_/X _15123_/Y _15094_/X _15123_/Y VGND VGND VPWR VPWR _15125_/B sky130_fd_sc_hd__a2bb2o_1
X_10597_ _10597_/A _09717_/X VGND VGND VPWR VPWR _10598_/A sky130_fd_sc_hd__or2b_1
X_12336_ _13397_/A _12336_/B VGND VGND VPWR VPWR _12336_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12267_ _12371_/A VGND VGND VPWR VPWR _12784_/A sky130_fd_sc_hd__buf_1
X_15055_ _15055_/A _15046_/X VGND VGND VPWR VPWR _15055_/X sky130_fd_sc_hd__or2b_1
X_14006_ _15418_/A _13959_/B _13959_/Y VGND VGND VPWR VPWR _14006_/Y sky130_fd_sc_hd__o21ai_1
X_11218_ _11085_/X _11217_/X _11085_/X _11217_/X VGND VGND VPWR VPWR _11219_/B sky130_fd_sc_hd__a2bb2o_1
X_12198_ _12198_/A _12251_/B VGND VGND VPWR VPWR _12198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11149_ _11148_/A _11147_/Y _11148_/Y _11147_/A _11529_/A VGND VGND VPWR VPWR _11316_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_95_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15957_ _15933_/X _15955_/X _16011_/B VGND VGND VPWR VPWR _15957_/X sky130_fd_sc_hd__o21a_1
X_15888_ _15888_/A _15888_/B VGND VGND VPWR VPWR _15888_/Y sky130_fd_sc_hd__nand2_1
X_14908_ _14908_/A _14908_/B VGND VGND VPWR VPWR _14908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14839_ _15051_/A _12372_/Y _12278_/Y _14752_/X VGND VGND VPWR VPWR _14839_/X sky130_fd_sc_hd__o22a_1
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08360_ input9/X _08279_/B _08359_/X VGND VGND VPWR VPWR _08361_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08291_ _08326_/A input33/X _08327_/A _08329_/A VGND VGND VPWR VPWR _08324_/A sky130_fd_sc_hd__o22a_1
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09814_ _09811_/X _08822_/A _09811_/X _08822_/A VGND VGND VPWR VPWR _09820_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09745_ _09745_/A _09745_/B VGND VGND VPWR VPWR _09791_/A sky130_fd_sc_hd__or2_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _13063_/A VGND VGND VPWR VPWR _11942_/A sky130_fd_sc_hd__buf_1
XFILLER_55_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _08650_/A _08627_/B VGND VGND VPWR VPWR _08634_/A sky130_fd_sc_hd__or2_1
XFILLER_27_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08558_ _08558_/A VGND VGND VPWR VPWR _08558_/Y sky130_fd_sc_hd__inv_2
X_08489_ _08336_/A _08260_/B _08475_/Y _08574_/A VGND VGND VPWR VPWR _08561_/A sky130_fd_sc_hd__o22a_1
X_10520_ _10906_/A _11595_/A VGND VGND VPWR VPWR _10625_/C sky130_fd_sc_hd__or2_1
X_10451_ _10448_/Y _12699_/A _10368_/X _10450_/Y VGND VGND VPWR VPWR _10451_/X sky130_fd_sc_hd__o22a_1
XFILLER_109_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13170_ _13106_/X _13169_/Y _13106_/X _13169_/Y VGND VGND VPWR VPWR _13188_/B sky130_fd_sc_hd__a2bb2o_1
X_10382_ _10370_/X _10381_/Y _10370_/X _10381_/Y VGND VGND VPWR VPWR _10450_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_124_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12121_ _13913_/A _12147_/B VGND VGND VPWR VPWR _12218_/A sky130_fd_sc_hd__and2_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12052_ _12042_/Y _12050_/X _12051_/Y VGND VGND VPWR VPWR _12052_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11003_ _11004_/A _11005_/B VGND VGND VPWR VPWR _11006_/A sky130_fd_sc_hd__and2_1
XFILLER_2_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15811_ _16110_/A _15811_/B VGND VGND VPWR VPWR _15811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15742_ _15678_/X _15741_/Y _15678_/X _15741_/Y VGND VGND VPWR VPWR _15811_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12954_ _12954_/A _12953_/X VGND VGND VPWR VPWR _12954_/X sky130_fd_sc_hd__or2b_1
XFILLER_58_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11905_ _11879_/Y _11903_/Y _11904_/Y VGND VGND VPWR VPWR _11906_/A sky130_fd_sc_hd__o21ai_1
X_15673_ _15673_/A _15673_/B VGND VGND VPWR VPWR _15673_/Y sky130_fd_sc_hd__nand2_1
X_12885_ _12938_/A VGND VGND VPWR VPWR _14476_/A sky130_fd_sc_hd__buf_1
XFILLER_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14580_/X _14623_/Y _14580_/X _14623_/Y VGND VGND VPWR VPWR _14653_/B sky130_fd_sc_hd__a2bb2o_1
X_11836_ _11836_/A _11836_/B VGND VGND VPWR VPWR _11836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _15261_/A VGND VGND VPWR VPWR _14577_/A sky130_fd_sc_hd__buf_1
X_11767_ _11767_/A _11767_/B VGND VGND VPWR VPWR _11768_/B sky130_fd_sc_hd__or2_1
XFILLER_14_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13506_ _13506_/A _13506_/B VGND VGND VPWR VPWR _13506_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10718_ _09651_/X _10717_/X _09651_/X _10717_/X VGND VGND VPWR VPWR _10719_/B sky130_fd_sc_hd__a2bb2oi_1
X_16225_ _16223_/A _16224_/A _16223_/Y _16224_/Y _16205_/A VGND VGND VPWR VPWR _16251_/A
+ sky130_fd_sc_hd__a221o_1
X_14486_ _14465_/X _14485_/Y _14465_/X _14485_/Y VGND VGND VPWR VPWR _14517_/B sky130_fd_sc_hd__a2bb2o_1
X_11698_ _13462_/A _11632_/B _11632_/Y _11636_/X VGND VGND VPWR VPWR _11698_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer2 _14275_/Y VGND VGND VPWR VPWR _14276_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13437_ _13437_/A _13437_/B VGND VGND VPWR VPWR _13437_/Y sky130_fd_sc_hd__nand2_1
X_10649_ _10584_/Y _10647_/Y _10648_/Y VGND VGND VPWR VPWR _10785_/A sky130_fd_sc_hd__o21ai_1
XFILLER_127_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16156_ _16113_/X _16155_/X _16113_/X _16155_/X VGND VGND VPWR VPWR _16157_/B sky130_fd_sc_hd__a2bb2oi_1
X_13368_ _13368_/A _13368_/B VGND VGND VPWR VPWR _13368_/X sky130_fd_sc_hd__or2_1
X_16087_ _16030_/A _16030_/B _16030_/Y VGND VGND VPWR VPWR _16087_/Y sky130_fd_sc_hd__o21ai_1
X_12319_ _12237_/X _12318_/Y _12237_/A _12318_/Y VGND VGND VPWR VPWR _12320_/B sky130_fd_sc_hd__a2bb2o_1
X_15107_ _15107_/A _15107_/B VGND VGND VPWR VPWR _15107_/Y sky130_fd_sc_hd__nand2_1
X_13299_ _13299_/A VGND VGND VPWR VPWR _13299_/Y sky130_fd_sc_hd__inv_2
X_15038_ _15038_/A _15038_/B VGND VGND VPWR VPWR _15038_/X sky130_fd_sc_hd__or2_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09530_ _09530_/A VGND VGND VPWR VPWR _09530_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09461_ _09459_/A _08639_/B _09459_/Y _09460_/Y VGND VGND VPWR VPWR _09461_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09392_ _09392_/A VGND VGND VPWR VPWR _09392_/X sky130_fd_sc_hd__clkbuf_2
X_08412_ _08717_/A VGND VGND VPWR VPWR _09251_/A sky130_fd_sc_hd__buf_1
XFILLER_24_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08343_ _08343_/A VGND VGND VPWR VPWR _08343_/Y sky130_fd_sc_hd__inv_2
X_08274_ input26/X VGND VGND VPWR VPWR _08275_/A sky130_fd_sc_hd__inv_4
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09728_ _09728_/A _09728_/B VGND VGND VPWR VPWR _09731_/B sky130_fd_sc_hd__or2_1
XFILLER_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09659_ _09597_/Y _09657_/X _09658_/Y VGND VGND VPWR VPWR _09659_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12670_ _10966_/Y _12669_/Y _10824_/Y VGND VGND VPWR VPWR _12671_/A sky130_fd_sc_hd__o21ai_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11623_/A VGND VGND VPWR VPWR _11621_/Y sky130_fd_sc_hd__inv_2
X_14340_ _14352_/A _14340_/B VGND VGND VPWR VPWR _15954_/A sky130_fd_sc_hd__or2_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11552_ _12396_/A _11652_/B VGND VGND VPWR VPWR _11552_/Y sky130_fd_sc_hd__nand2_1
X_14271_ _15860_/A _14271_/B VGND VGND VPWR VPWR _14271_/Y sky130_fd_sc_hd__nand2_1
X_11483_ _14744_/A _11482_/B _11482_/X _11280_/X VGND VGND VPWR VPWR _11483_/X sky130_fd_sc_hd__o22a_1
X_10503_ _11783_/A _10409_/B _11783_/A _10409_/B VGND VGND VPWR VPWR _10503_/X sky130_fd_sc_hd__a2bb2o_1
X_16010_ _16040_/A _16040_/B VGND VGND VPWR VPWR _16010_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13222_ _14673_/A VGND VGND VPWR VPWR _14740_/A sky130_fd_sc_hd__buf_1
X_10434_ _13563_/A _10400_/B _10400_/X _10433_/X VGND VGND VPWR VPWR _10434_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13153_ _13200_/A _13200_/B VGND VGND VPWR VPWR _13153_/Y sky130_fd_sc_hd__nor2_1
X_10365_ _10367_/A VGND VGND VPWR VPWR _10365_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12104_ _12103_/A _12160_/B _12103_/Y VGND VGND VPWR VPWR _12104_/Y sky130_fd_sc_hd__o21ai_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ _13760_/A VGND VGND VPWR VPWR _15261_/A sky130_fd_sc_hd__buf_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10296_/A VGND VGND VPWR VPWR _10325_/A sky130_fd_sc_hd__inv_2
X_12035_ _11969_/X _12034_/Y _11969_/X _12034_/Y VGND VGND VPWR VPWR _12055_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13986_ _13861_/X _13883_/A _13882_/X VGND VGND VPWR VPWR _13986_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15725_ _15817_/A _15817_/B VGND VGND VPWR VPWR _15725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12937_ _12892_/Y _12935_/X _12936_/Y VGND VGND VPWR VPWR _12937_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15656_ _15656_/A VGND VGND VPWR VPWR _16028_/A sky130_fd_sc_hd__clkinvlp_2
X_12868_ _12948_/A _12949_/B VGND VGND VPWR VPWR _12868_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14607_ _14664_/A _14664_/B _14606_/Y VGND VGND VPWR VPWR _14607_/Y sky130_fd_sc_hd__o21ai_1
X_11819_ _10440_/A _11848_/B _10440_/A _11848_/B VGND VGND VPWR VPWR _11819_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15587_ _15545_/X _15586_/X _15545_/X _15586_/X VGND VGND VPWR VPWR _15588_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12857_/A _12857_/B VGND VGND VPWR VPWR _12799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14538_ _14587_/A _14587_/B VGND VGND VPWR VPWR _14538_/Y sky130_fd_sc_hd__nor2_1
X_14469_ _14441_/Y _14467_/X _14468_/Y VGND VGND VPWR VPWR _14469_/X sky130_fd_sc_hd__o21a_1
X_16208_ _16208_/A VGND VGND VPWR VPWR _16208_/Y sky130_fd_sc_hd__inv_2
X_16139_ _16139_/A VGND VGND VPWR VPWR _16139_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08961_ _08957_/Y _11399_/A _08960_/Y VGND VGND VPWR VPWR _08968_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08892_ _08686_/X _08891_/X _08686_/X _08891_/X VGND VGND VPWR VPWR _08976_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09513_ _09490_/A _09490_/B _09490_/Y _09512_/X VGND VGND VPWR VPWR _09513_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09444_ _10907_/A VGND VGND VPWR VPWR _09445_/A sky130_fd_sc_hd__clkbuf_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09375_ _10239_/A VGND VGND VPWR VPWR _09376_/B sky130_fd_sc_hd__buf_1
X_08326_ _08326_/A input33/X VGND VGND VPWR VPWR _08327_/B sky130_fd_sc_hd__nor2_1
X_08257_ input16/X _08257_/B VGND VGND VPWR VPWR _08332_/A sky130_fd_sc_hd__nor2_1
XFILLER_125_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10150_ _08786_/B _10130_/B _10131_/B VGND VGND VPWR VPWR _10151_/B sky130_fd_sc_hd__a21bo_1
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10081_ _10081_/A _10081_/B VGND VGND VPWR VPWR _10969_/B sky130_fd_sc_hd__or2_1
XFILLER_102_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13840_ _13831_/Y _13838_/X _13839_/Y VGND VGND VPWR VPWR _13840_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13771_ _13806_/A _13769_/X _13770_/X VGND VGND VPWR VPWR _13771_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10983_ _10983_/A _10983_/B VGND VGND VPWR VPWR _10983_/Y sky130_fd_sc_hd__nand2_1
X_15510_ _15510_/A VGND VGND VPWR VPWR _15510_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12722_ _12681_/X _12721_/X _12681_/X _12721_/X VGND VGND VPWR VPWR _13457_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15441_ _15441_/A _15416_/X VGND VGND VPWR VPWR _15441_/X sky130_fd_sc_hd__or2b_1
XFILLER_43_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12653_ _15285_/A VGND VGND VPWR VPWR _13984_/A sky130_fd_sc_hd__inv_2
X_12584_ _12581_/Y _12583_/Y _12581_/A _12583_/A _12502_/A VGND VGND VPWR VPWR _12622_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_90_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15372_ _15372_/A _15343_/X VGND VGND VPWR VPWR _15372_/X sky130_fd_sc_hd__or2b_1
X_11604_ _11619_/A VGND VGND VPWR VPWR _12680_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14323_ _15960_/A _14389_/B VGND VGND VPWR VPWR _14323_/X sky130_fd_sc_hd__and2_1
X_11535_ _09370_/B _10238_/B _10238_/X VGND VGND VPWR VPWR _11536_/B sky130_fd_sc_hd__a21boi_1
XFILLER_7_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14254_ _14227_/Y _14252_/Y _14253_/Y VGND VGND VPWR VPWR _14255_/A sky130_fd_sc_hd__o21ai_2
XFILLER_7_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11466_ _14143_/A VGND VGND VPWR VPWR _13447_/A sky130_fd_sc_hd__buf_1
X_13205_ _13147_/Y _13203_/X _13204_/Y VGND VGND VPWR VPWR _13205_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14185_ _15857_/A _14274_/B VGND VGND VPWR VPWR _14185_/Y sky130_fd_sc_hd__nor2_1
X_10417_ _10517_/A VGND VGND VPWR VPWR _12827_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11397_ _11397_/A VGND VGND VPWR VPWR _11397_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13136_ _13139_/A VGND VGND VPWR VPWR _15289_/A sky130_fd_sc_hd__buf_1
X_10348_ _10454_/A _11714_/B VGND VGND VPWR VPWR _10349_/A sky130_fd_sc_hd__nand2_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13067_ _15249_/A _13115_/B VGND VGND VPWR VPWR _13067_/Y sky130_fd_sc_hd__nor2_1
X_10279_ _11716_/A VGND VGND VPWR VPWR _11723_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_3_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12018_ _11942_/A _11978_/B _11978_/Y VGND VGND VPWR VPWR _12018_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13969_ _13873_/A _13868_/X _13873_/B VGND VGND VPWR VPWR _13969_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_53_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15708_ _14927_/X _15707_/X _14927_/X _15707_/X VGND VGND VPWR VPWR _15709_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_80_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15639_ _15639_/A _15519_/X VGND VGND VPWR VPWR _15641_/A sky130_fd_sc_hd__or2b_1
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09160_ _09160_/A VGND VGND VPWR VPWR _09160_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09091_ _10016_/B _09073_/B _09074_/B VGND VGND VPWR VPWR _09703_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09993_ _09993_/A _09993_/B VGND VGND VPWR VPWR _09993_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08944_ _08944_/A _08944_/B VGND VGND VPWR VPWR _08944_/X sky130_fd_sc_hd__or2_1
XFILLER_111_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08875_ _08984_/A _08984_/B VGND VGND VPWR VPWR _08875_/X sky130_fd_sc_hd__and2_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09427_ _09426_/A _09433_/B _09426_/Y VGND VGND VPWR VPWR _09428_/A sky130_fd_sc_hd__o21ai_1
XFILLER_100_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09358_ _09478_/B _09863_/A _09346_/Y _09357_/X VGND VGND VPWR VPWR _09358_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08309_ _08309_/A VGND VGND VPWR VPWR _08309_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11320_ _11607_/A _11320_/B VGND VGND VPWR VPWR _11321_/A sky130_fd_sc_hd__or2_1
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09289_ _08922_/B _08936_/Y _08922_/B _08936_/Y VGND VGND VPWR VPWR _10230_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11251_ _11413_/A _11251_/B _13935_/B VGND VGND VPWR VPWR _11251_/X sky130_fd_sc_hd__or3_1
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10202_ _09403_/X _08931_/Y _09404_/Y _08931_/A VGND VGND VPWR VPWR _11245_/A sky130_fd_sc_hd__a22o_2
X_11182_ _09140_/Y _11181_/A _09140_/A _11181_/Y _09204_/X VGND VGND VPWR VPWR _13366_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_133_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10133_ _10133_/A _10133_/B VGND VGND VPWR VPWR _10134_/B sky130_fd_sc_hd__or2_1
XFILLER_121_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15990_ _15991_/A _15991_/B VGND VGND VPWR VPWR _15990_/X sky130_fd_sc_hd__and2_1
XFILLER_95_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14941_ _14939_/Y _14940_/X _14939_/Y _14940_/X VGND VGND VPWR VPWR _14980_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10064_ _10063_/A _10063_/B _09963_/A _10063_/X VGND VGND VPWR VPWR _10067_/A sky130_fd_sc_hd__a22o_1
X_14872_ _14872_/A VGND VGND VPWR VPWR _15546_/A sky130_fd_sc_hd__buf_1
XFILLER_90_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13823_ _14630_/A _13843_/B VGND VGND VPWR VPWR _13823_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13754_ _13754_/A VGND VGND VPWR VPWR _13754_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10966_ _12084_/A _10966_/B VGND VGND VPWR VPWR _10966_/Y sky130_fd_sc_hd__nor2_1
X_16473_ _16473_/D _16454_/Y VGND VGND VPWR VPWR _16473_/Q sky130_fd_sc_hd__dlxtn_1
X_13685_ _13685_/A VGND VGND VPWR VPWR _13685_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12705_ _12705_/A VGND VGND VPWR VPWR _12705_/Y sky130_fd_sc_hd__inv_2
X_10897_ _09296_/A _10896_/A _09296_/Y _10896_/Y _09445_/A VGND VGND VPWR VPWR _13828_/A
+ sky130_fd_sc_hd__a221o_4
X_12636_ _12636_/A _12636_/B VGND VGND VPWR VPWR _12636_/X sky130_fd_sc_hd__or2_1
X_15424_ _15286_/X _15423_/X _15286_/X _15423_/X VGND VGND VPWR VPWR _15424_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15355_ _15290_/X _15354_/X _15290_/X _15354_/X VGND VGND VPWR VPWR _15422_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12567_ _15529_/A VGND VGND VPWR VPWR _14912_/A sky130_fd_sc_hd__buf_1
X_14306_ _13441_/A _13441_/B _13441_/Y VGND VGND VPWR VPWR _14306_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12498_ _12491_/X _12497_/X _12491_/X _12497_/X VGND VGND VPWR VPWR _12498_/X sky130_fd_sc_hd__a2bb2o_1
X_15286_ _15287_/A _15284_/Y _15287_/B VGND VGND VPWR VPWR _15286_/X sky130_fd_sc_hd__o21ba_1
X_11518_ _12376_/A VGND VGND VPWR VPWR _12275_/A sky130_fd_sc_hd__inv_2
XFILLER_8_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14237_ _15509_/A _14081_/B _14081_/Y VGND VGND VPWR VPWR _14238_/A sky130_fd_sc_hd__a21oi_1
XFILLER_109_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11449_ _15534_/A _11449_/B VGND VGND VPWR VPWR _11449_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14168_ _14139_/X _14167_/Y _14139_/X _14167_/Y VGND VGND VPWR VPWR _14169_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_98_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13119_ _15243_/A _13119_/B VGND VGND VPWR VPWR _13119_/Y sky130_fd_sc_hd__nand2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14051_/X _14098_/X _14051_/X _14098_/X VGND VGND VPWR VPWR _14099_/Y sky130_fd_sc_hd__a2bb2oi_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08660_ _08660_/A _08662_/B VGND VGND VPWR VPWR _08919_/A sky130_fd_sc_hd__or2b_1
XFILLER_94_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08591_ _08794_/A _09213_/B _08794_/A _09213_/B VGND VGND VPWR VPWR _08592_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09212_ _09212_/A VGND VGND VPWR VPWR _09212_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09143_ _09432_/A _09175_/B VGND VGND VPWR VPWR _09143_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09074_ _10015_/B _09074_/B VGND VGND VPWR VPWR _09075_/B sky130_fd_sc_hd__or2_1
XFILLER_116_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09976_ _09971_/Y _09974_/Y _09975_/Y VGND VGND VPWR VPWR _09978_/B sky130_fd_sc_hd__o21ai_1
X_08927_ _10102_/A _09680_/A VGND VGND VPWR VPWR _08928_/A sky130_fd_sc_hd__or2_2
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08858_ _09502_/A _08842_/Y _08844_/Y _08857_/X VGND VGND VPWR VPWR _08955_/A sky130_fd_sc_hd__o22a_1
XFILLER_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08789_ _08789_/A VGND VGND VPWR VPWR _08789_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10820_ _10242_/B _10155_/B _10155_/Y VGND VGND VPWR VPWR _10821_/A sky130_fd_sc_hd__a21oi_1
XFILLER_13_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10751_ _10751_/A VGND VGND VPWR VPWR _10751_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13470_ _13458_/X _13469_/X _13458_/X _13469_/X VGND VGND VPWR VPWR _13470_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_13_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12421_ _12683_/A _12420_/B _12420_/X _12382_/B VGND VGND VPWR VPWR _12422_/B sky130_fd_sc_hd__a22o_1
X_10682_ _10682_/A VGND VGND VPWR VPWR _11994_/A sky130_fd_sc_hd__inv_2
X_12352_ _12348_/Y _12551_/A _12351_/Y VGND VGND VPWR VPWR _12543_/A sky130_fd_sc_hd__o21ai_2
X_15140_ _15140_/A _15140_/B VGND VGND VPWR VPWR _15140_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11303_ _13780_/A VGND VGND VPWR VPWR _13788_/A sky130_fd_sc_hd__buf_1
X_12283_ _13788_/A _12367_/B VGND VGND VPWR VPWR _12283_/Y sky130_fd_sc_hd__nand2_1
X_15071_ _15035_/X _15070_/X _15035_/X _15070_/X VGND VGND VPWR VPWR _15072_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11234_ _12229_/A VGND VGND VPWR VPWR _14038_/A sky130_fd_sc_hd__buf_1
X_14022_ _13948_/X _14021_/Y _13948_/X _14021_/Y VGND VGND VPWR VPWR _14023_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11165_ _13715_/A _11297_/B _11164_/Y VGND VGND VPWR VPWR _11165_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15973_ _15915_/X _15971_/X _15993_/B VGND VGND VPWR VPWR _15973_/X sky130_fd_sc_hd__o21a_1
X_11096_ _09432_/B _09382_/B _09382_/X VGND VGND VPWR VPWR _11097_/B sky130_fd_sc_hd__a21boi_1
X_10116_ _10116_/A _10116_/B VGND VGND VPWR VPWR _10117_/A sky130_fd_sc_hd__or2_1
X_14924_ _15548_/A _14924_/B VGND VGND VPWR VPWR _14924_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10047_ _10047_/A _10047_/B VGND VGND VPWR VPWR _10047_/Y sky130_fd_sc_hd__nor2_1
X_14855_ _15353_/A _14958_/B _14854_/Y VGND VGND VPWR VPWR _14855_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08231__2 _16357_/A VGND VGND VPWR VPWR _08232_/A sky130_fd_sc_hd__inv_2
X_14786_ _14786_/A _14786_/B VGND VGND VPWR VPWR _14786_/X sky130_fd_sc_hd__and2_1
XFILLER_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13806_ _13806_/A _13770_/X VGND VGND VPWR VPWR _13806_/X sky130_fd_sc_hd__or2b_1
X_11998_ _11999_/A _11999_/B VGND VGND VPWR VPWR _11998_/X sky130_fd_sc_hd__and2_1
X_13737_ _13764_/A _13764_/B VGND VGND VPWR VPWR _13815_/A sky130_fd_sc_hd__and2_1
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10949_ _10949_/A _10949_/B VGND VGND VPWR VPWR _10949_/Y sky130_fd_sc_hd__nor2_1
X_16456_ VGND VGND VPWR VPWR _16456_/HI _16456_/LO sky130_fd_sc_hd__conb_1
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15407_ _15456_/A _15405_/X _15406_/X VGND VGND VPWR VPWR _15407_/X sky130_fd_sc_hd__o21a_1
X_13668_ _13623_/A _13667_/Y _13623_/A _13667_/Y VGND VGND VPWR VPWR _13692_/B sky130_fd_sc_hd__a2bb2o_1
X_16387_ _16124_/X _16386_/X _16124_/X _16386_/X VGND VGND VPWR VPWR _16388_/B sky130_fd_sc_hd__a2bb2o_1
X_12619_ _14231_/A _14235_/A _12618_/X VGND VGND VPWR VPWR _12619_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13599_ _13563_/A _13563_/B _13564_/A VGND VGND VPWR VPWR _13599_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_117_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15338_ _15381_/A _15336_/X _15337_/X VGND VGND VPWR VPWR _15338_/X sky130_fd_sc_hd__o21a_1
XANTENNA_0 _16472_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15269_ _15212_/X _15268_/X _15212_/X _15268_/X VGND VGND VPWR VPWR _15270_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _09830_/A VGND VGND VPWR VPWR _09830_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09736_/A _09736_/B _09739_/A VGND VGND VPWR VPWR _10046_/A sky130_fd_sc_hd__a21bo_1
XFILLER_39_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08712_/A _09470_/B VGND VGND VPWR VPWR _08712_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09692_ _09692_/A _09692_/B VGND VGND VPWR VPWR _09695_/A sky130_fd_sc_hd__or2_1
Xrebuffer12 rebuffer13/X VGND VGND VPWR VPWR rebuffer12/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08643_ _08718_/A VGND VGND VPWR VPWR _09458_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer45 _10001_/B1 VGND VGND VPWR VPWR _11599_/B1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer34 _10190_/X VGND VGND VPWR VPWR _11324_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer23 _10191_/X VGND VGND VPWR VPWR _11528_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer56 _10283_/B2 VGND VGND VPWR VPWR _12708_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_35_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08574_ _08574_/A VGND VGND VPWR VPWR _08574_/Y sky130_fd_sc_hd__clkinvlp_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09126_ _09701_/A _09126_/B VGND VGND VPWR VPWR _09126_/Y sky130_fd_sc_hd__nand2_1
X_09057_ _08789_/Y _09050_/A _08789_/A _09050_/Y VGND VGND VPWR VPWR _10013_/B sky130_fd_sc_hd__o22a_1
XFILLER_116_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09959_ _09951_/Y _09957_/Y _09958_/Y VGND VGND VPWR VPWR _09972_/B sky130_fd_sc_hd__o21ai_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12970_ _12941_/X _12969_/Y _12941_/X _12969_/Y VGND VGND VPWR VPWR _13029_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11921_ _11921_/A _11921_/B VGND VGND VPWR VPWR _11921_/X sky130_fd_sc_hd__or2_1
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14640_ _14645_/A _14645_/B VGND VGND VPWR VPWR _14715_/A sky130_fd_sc_hd__and2_1
X_11852_ _11850_/A _11850_/B _11850_/X _11851_/Y VGND VGND VPWR VPWR _11916_/B sky130_fd_sc_hd__a22o_1
X_14571_ _15270_/A _14571_/B VGND VGND VPWR VPWR _14571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10803_ _10953_/A VGND VGND VPWR VPWR _11009_/A sky130_fd_sc_hd__buf_1
XFILLER_26_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16310_ _16250_/X _16309_/Y _16250_/X _16309_/Y VGND VGND VPWR VPWR _16318_/B sky130_fd_sc_hd__o2bb2a_1
X_11783_ _11783_/A _11783_/B VGND VGND VPWR VPWR _11783_/X sky130_fd_sc_hd__and2_1
X_13522_ _13524_/A VGND VGND VPWR VPWR _15032_/A sky130_fd_sc_hd__buf_1
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10734_ _09960_/A _09645_/B _09645_/Y VGND VGND VPWR VPWR _10736_/A sky130_fd_sc_hd__o21ai_1
X_16241_ _16241_/A VGND VGND VPWR VPWR _16241_/Y sky130_fd_sc_hd__clkinvlp_2
X_13453_ _13450_/X _13452_/Y _13450_/X _13452_/Y VGND VGND VPWR VPWR _13453_/X sky130_fd_sc_hd__a2bb2o_1
X_10665_ _10664_/A _10664_/B _10664_/Y _09392_/A VGND VGND VPWR VPWR _11016_/A sky130_fd_sc_hd__o211a_1
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16172_ _16109_/X _16171_/X _16109_/X _16171_/X VGND VGND VPWR VPWR _16173_/B sky130_fd_sc_hd__a2bb2oi_1
X_13384_ _13384_/A _13366_/X VGND VGND VPWR VPWR _13384_/X sky130_fd_sc_hd__or2b_1
X_12404_ _13544_/A _12404_/B VGND VGND VPWR VPWR _12405_/B sky130_fd_sc_hd__or2_1
XFILLER_127_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12335_ _12241_/X _12334_/Y _12241_/X _12334_/Y VGND VGND VPWR VPWR _12581_/A sky130_fd_sc_hd__a2bb2o_1
X_10596_ _11904_/A _10642_/B VGND VGND VPWR VPWR _10596_/Y sky130_fd_sc_hd__nor2_1
X_15123_ _15066_/A _15066_/B _15066_/Y VGND VGND VPWR VPWR _15123_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15054_ _15054_/A _15054_/B VGND VGND VPWR VPWR _15054_/Y sky130_fd_sc_hd__nand2_1
X_12266_ _13500_/A VGND VGND VPWR VPWR _12371_/A sky130_fd_sc_hd__inv_2
X_14005_ _14005_/A _14065_/B VGND VGND VPWR VPWR _14140_/A sky130_fd_sc_hd__and2_1
X_11217_ _11217_/A _11086_/X VGND VGND VPWR VPWR _11217_/X sky130_fd_sc_hd__or2b_1
X_12197_ _12161_/X _12196_/Y _12161_/X _12196_/Y VGND VGND VPWR VPWR _12251_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11148_ _11148_/A VGND VGND VPWR VPWR _11148_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15956_ _15956_/A _15956_/B VGND VGND VPWR VPWR _16011_/B sky130_fd_sc_hd__or2_1
X_11079_ _11242_/A _11076_/X _11078_/X VGND VGND VPWR VPWR _11079_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15887_ _15883_/Y _15885_/X _15886_/Y VGND VGND VPWR VPWR _15887_/X sky130_fd_sc_hd__o21a_1
X_14907_ _14901_/Y _14905_/X _14906_/Y VGND VGND VPWR VPWR _14907_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14838_ _14754_/A _14754_/B _14751_/X _14754_/Y VGND VGND VPWR VPWR _14838_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14769_ _14743_/X _14768_/Y _14743_/X _14768_/Y VGND VGND VPWR VPWR _14771_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08290_ _08331_/A input32/X _08332_/A _08334_/A VGND VGND VPWR VPWR _08329_/A sky130_fd_sc_hd__o22a_1
XFILLER_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16439_ _16419_/B _16436_/X _16435_/X _16438_/X VGND VGND VPWR VPWR _16439_/X sky130_fd_sc_hd__o22a_1
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09813_ _09812_/X _08813_/A _09812_/X _08813_/A VGND VGND VPWR VPWR _09821_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09744_ _08524_/Y _09743_/X _08524_/Y _09743_/X VGND VGND VPWR VPWR _09745_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09675_ _10933_/A _09675_/B VGND VGND VPWR VPWR _13063_/A sky130_fd_sc_hd__or2_2
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _08625_/A _08365_/Y _08625_/Y _08365_/A VGND VGND VPWR VPWR _08627_/B sky130_fd_sc_hd__o22a_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08557_ _09737_/A _08567_/B VGND VGND VPWR VPWR _08558_/A sky130_fd_sc_hd__or2_1
XFILLER_52_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08488_ _08263_/A _08341_/B _08476_/Y _08587_/A VGND VGND VPWR VPWR _08574_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10450_ _10450_/A _11767_/A VGND VGND VPWR VPWR _10450_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09109_ _09714_/A _09107_/B _09107_/X _09108_/Y VGND VGND VPWR VPWR _09113_/B sky130_fd_sc_hd__o22ai_2
X_10381_ _10381_/A VGND VGND VPWR VPWR _10381_/Y sky130_fd_sc_hd__clkinvlp_2
X_12120_ _12058_/X _12119_/Y _12058_/X _12119_/Y VGND VGND VPWR VPWR _12147_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12051_ _13828_/A _12051_/B VGND VGND VPWR VPWR _12051_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11002_ _10932_/X _11001_/Y _10932_/X _11001_/Y VGND VGND VPWR VPWR _11005_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15810_ _15749_/Y _15808_/X _15809_/Y VGND VGND VPWR VPWR _15810_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15741_ _15679_/A _15679_/B _15679_/Y VGND VGND VPWR VPWR _15741_/Y sky130_fd_sc_hd__o21ai_1
X_12953_ _14948_/A _12953_/B VGND VGND VPWR VPWR _12953_/X sky130_fd_sc_hd__or2_1
X_15672_ _15638_/Y _15670_/X _15671_/Y VGND VGND VPWR VPWR _15672_/X sky130_fd_sc_hd__o21a_1
XFILLER_73_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11904_ _11904_/A _11904_/B VGND VGND VPWR VPWR _11904_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14623_ _14581_/A _14581_/B _14581_/Y VGND VGND VPWR VPWR _14623_/Y sky130_fd_sc_hd__o21ai_1
X_12884_ _14531_/A _12940_/B VGND VGND VPWR VPWR _12884_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11795_/X _11834_/X _11795_/X _11834_/X VGND VGND VPWR VPWR _11836_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14579_/A _14579_/B VGND VGND VPWR VPWR _14554_/Y sky130_fd_sc_hd__nor2_1
X_11766_ _11767_/A _11767_/B VGND VGND VPWR VPWR _11766_/X sky130_fd_sc_hd__and2_1
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _14466_/A _14466_/B _14466_/Y VGND VGND VPWR VPWR _14485_/Y sky130_fd_sc_hd__o21ai_1
X_13505_ _10988_/X _13488_/X _10988_/X _13488_/X VGND VGND VPWR VPWR _13506_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10717_ _09978_/A _09652_/B _09652_/Y VGND VGND VPWR VPWR _10717_/X sky130_fd_sc_hd__o21a_1
X_16224_ _16224_/A VGND VGND VPWR VPWR _16224_/Y sky130_fd_sc_hd__inv_2
X_13436_ _13432_/Y _13434_/Y _13435_/Y VGND VGND VPWR VPWR _13436_/X sky130_fd_sc_hd__o21a_1
X_11697_ _13994_/A VGND VGND VPWR VPWR _13462_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10648_ _11910_/A _10648_/B VGND VGND VPWR VPWR _10648_/Y sky130_fd_sc_hd__nand2_1
Xrebuffer3 rebuffer4/X VGND VGND VPWR VPWR rebuffer3/X sky130_fd_sc_hd__dlygate4sd1_1
X_16155_ _16067_/X _16155_/B VGND VGND VPWR VPWR _16155_/X sky130_fd_sc_hd__and2b_1
X_13367_ _13384_/A _13365_/X _13366_/X VGND VGND VPWR VPWR _13367_/X sky130_fd_sc_hd__o21a_1
X_10579_ _10545_/X _10661_/B _10545_/X _10661_/B VGND VGND VPWR VPWR _10579_/X sky130_fd_sc_hd__a2bb2o_1
X_16086_ _16086_/A _16089_/B VGND VGND VPWR VPWR _16086_/Y sky130_fd_sc_hd__nor2_1
X_12318_ _13350_/A _12238_/B _12238_/Y VGND VGND VPWR VPWR _12318_/Y sky130_fd_sc_hd__o21ai_1
X_13298_ _13230_/Y _13296_/Y _13297_/Y VGND VGND VPWR VPWR _13299_/A sky130_fd_sc_hd__o21ai_1
X_15106_ _15100_/X _15105_/Y _15100_/X _15105_/Y VGND VGND VPWR VPWR _15107_/B sky130_fd_sc_hd__a2bb2o_1
X_12249_ _14061_/A _12205_/B _12205_/Y _12248_/X VGND VGND VPWR VPWR _12249_/X sky130_fd_sc_hd__a2bb2o_1
X_15037_ _15070_/A _15035_/X _15036_/X VGND VGND VPWR VPWR _15037_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15939_ _15952_/A _15952_/B VGND VGND VPWR VPWR _15939_/X sky130_fd_sc_hd__and2_1
XFILLER_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09460_ _09460_/A VGND VGND VPWR VPWR _09460_/Y sky130_fd_sc_hd__inv_2
X_08411_ _09225_/A VGND VGND VPWR VPWR _08717_/A sky130_fd_sc_hd__inv_2
XFILLER_24_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09391_ _09391_/A VGND VGND VPWR VPWR _09392_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08342_ _08342_/A _08342_/B VGND VGND VPWR VPWR _08343_/A sky130_fd_sc_hd__or2_1
X_08273_ input10/X VGND VGND VPWR VPWR _08357_/B sky130_fd_sc_hd__inv_2
XFILLER_20_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09727_ _09727_/A VGND VGND VPWR VPWR _09727_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09658_ _09987_/A _09658_/B VGND VGND VPWR VPWR _09658_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _16357_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08609_ _08609_/A VGND VGND VPWR VPWR _10113_/B sky130_fd_sc_hd__inv_2
X_09589_ _08688_/A _09019_/A _09532_/A VGND VGND VPWR VPWR _09589_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _12680_/A _11619_/B _11619_/Y VGND VGND VPWR VPWR _11620_/Y sky130_fd_sc_hd__a21oi_1
X_11551_ _11495_/X _11550_/Y _11495_/X _11550_/Y VGND VGND VPWR VPWR _11652_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10502_ _11840_/A VGND VGND VPWR VPWR _13605_/A sky130_fd_sc_hd__buf_1
X_14270_ _14270_/A VGND VGND VPWR VPWR _14270_/Y sky130_fd_sc_hd__inv_2
X_11482_ _11482_/A _11482_/B VGND VGND VPWR VPWR _11482_/X sky130_fd_sc_hd__and2_1
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13221_ _15057_/A VGND VGND VPWR VPWR _14673_/A sky130_fd_sc_hd__inv_2
X_10433_ _13567_/A _10409_/B _10409_/X _10432_/X VGND VGND VPWR VPWR _10433_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13152_ _13118_/X _13151_/Y _13118_/X _13151_/Y VGND VGND VPWR VPWR _13200_/B sky130_fd_sc_hd__a2bb2o_1
X_10364_ _11758_/A VGND VGND VPWR VPWR _13521_/A sky130_fd_sc_hd__buf_1
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12103_ _12103_/A _12160_/B VGND VGND VPWR VPWR _12103_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13083_ _13083_/A VGND VGND VPWR VPWR _13760_/A sky130_fd_sc_hd__inv_2
X_10295_ _12707_/A _10291_/B _10291_/X _10294_/Y VGND VGND VPWR VPWR _10295_/X sky130_fd_sc_hd__a22o_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12034_ _13083_/A _11970_/B _11970_/Y VGND VGND VPWR VPWR _12034_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13985_ _13983_/X _13985_/B VGND VGND VPWR VPWR _13985_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15724_ _15684_/X _15723_/Y _15684_/X _15723_/Y VGND VGND VPWR VPWR _15817_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12936_ _12936_/A _12936_/B VGND VGND VPWR VPWR _12936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15655_ _15781_/A _15655_/B VGND VGND VPWR VPWR _15656_/A sky130_fd_sc_hd__or2_1
X_12867_ _12860_/X _12866_/Y _12860_/X _12866_/Y VGND VGND VPWR VPWR _12949_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15586_ _15500_/X _15586_/B VGND VGND VPWR VPWR _15586_/X sky130_fd_sc_hd__and2b_1
X_14606_ _14664_/A _14664_/B VGND VGND VPWR VPWR _14606_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11818_ _11850_/B _11817_/Y _11850_/B _11817_/Y VGND VGND VPWR VPWR _11848_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14522_/X _14536_/X _14522_/X _14536_/X VGND VGND VPWR VPWR _14587_/B sky130_fd_sc_hd__a2bb2o_1
X_12798_ _12781_/X _12797_/Y _12781_/X _12797_/Y VGND VGND VPWR VPWR _12857_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11749_ _11748_/A _11748_/B _10224_/B _11748_/X VGND VGND VPWR VPWR _11750_/A sky130_fd_sc_hd__a22o_1
X_14468_ _14468_/A _14468_/B VGND VGND VPWR VPWR _14468_/Y sky130_fd_sc_hd__nand2_1
X_16207_ _16207_/A VGND VGND VPWR VPWR _16207_/Y sky130_fd_sc_hd__inv_2
X_14399_ _14284_/X _14398_/Y _14284_/X _14398_/Y VGND VGND VPWR VPWR _14399_/Y sky130_fd_sc_hd__a2bb2oi_1
X_13419_ _13357_/X _13418_/X _13357_/X _13418_/X VGND VGND VPWR VPWR _13419_/Y sky130_fd_sc_hd__a2bb2oi_1
X_16138_ _16138_/A _16121_/X VGND VGND VPWR VPWR _16139_/A sky130_fd_sc_hd__or2b_1
XFILLER_130_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16069_ _16043_/X _16068_/Y _16043_/X _16068_/Y VGND VGND VPWR VPWR _16112_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08960_ _08960_/A _08960_/B VGND VGND VPWR VPWR _08960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08891_ _09555_/A _08571_/A _08573_/A VGND VGND VPWR VPWR _08891_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09512_ _08795_/X _09492_/B _09492_/Y _09511_/X VGND VGND VPWR VPWR _09512_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09443_ _09441_/X _09442_/X _09441_/X _09442_/X VGND VGND VPWR VPWR _10907_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_24_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09374_ _09335_/X _08878_/Y _09335_/X _08878_/Y VGND VGND VPWR VPWR _10239_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08325_ _08323_/Y _08324_/A _08323_/A _08324_/Y _08304_/X VGND VGND VPWR VPWR _08555_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08256_ input32/X VGND VGND VPWR VPWR _08257_/B sky130_fd_sc_hd__inv_2
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10080_ _10049_/X _10078_/X _10816_/B VGND VGND VPWR VPWR _10080_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13770_ _13770_/A _13770_/B VGND VGND VPWR VPWR _13770_/X sky130_fd_sc_hd__or2_1
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10982_ _09327_/B _10241_/B _10241_/X VGND VGND VPWR VPWR _10983_/B sky130_fd_sc_hd__a21boi_1
X_12721_ _12683_/A _12683_/B _12683_/Y _12720_/X VGND VGND VPWR VPWR _12721_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12652_ _12642_/Y _12650_/Y _14162_/B VGND VGND VPWR VPWR _12652_/Y sky130_fd_sc_hd__o21ai_1
X_15440_ _15440_/A _15440_/B VGND VGND VPWR VPWR _15440_/X sky130_fd_sc_hd__and2_1
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11603_ _11602_/A _11602_/B _11602_/Y _10984_/X VGND VGND VPWR VPWR _11619_/A sky130_fd_sc_hd__o211a_1
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12583_ _12583_/A VGND VGND VPWR VPWR _12583_/Y sky130_fd_sc_hd__inv_2
X_15371_ _15412_/A _15412_/B VGND VGND VPWR VPWR _15447_/A sky130_fd_sc_hd__and2_1
XFILLER_11_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14322_ _14267_/A _14321_/Y _14267_/A _14321_/Y VGND VGND VPWR VPWR _14389_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11534_ _11522_/X _11533_/Y _11522_/X _11533_/Y VGND VGND VPWR VPWR _11623_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14253_ _15878_/A _14253_/B VGND VGND VPWR VPWR _14253_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11465_ _12410_/A VGND VGND VPWR VPWR _14143_/A sky130_fd_sc_hd__buf_1
XFILLER_7_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13204_ _13204_/A _13204_/B VGND VGND VPWR VPWR _13204_/Y sky130_fd_sc_hd__nand2_1
X_10416_ _08402_/X _10277_/A _08929_/A _10339_/Y _10420_/B VGND VGND VPWR VPWR _10517_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14184_ _12633_/X _14183_/X _12633_/X _14183_/X VGND VGND VPWR VPWR _14274_/B sky130_fd_sc_hd__a2bb2o_1
X_11396_ _08968_/A _08968_/B _08968_/Y VGND VGND VPWR VPWR _11397_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13135_ _15167_/A VGND VGND VPWR VPWR _14934_/A sky130_fd_sc_hd__clkbuf_2
X_10347_ _10347_/A VGND VGND VPWR VPWR _11714_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13066_ _13024_/X _13065_/X _13024_/X _13065_/X VGND VGND VPWR VPWR _13115_/B sky130_fd_sc_hd__a2bb2o_1
X_10278_ _08929_/A _10277_/A _08402_/X _10277_/Y _10268_/A VGND VGND VPWR VPWR _11716_/A
+ sky130_fd_sc_hd__o221a_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12017_ _12063_/A VGND VGND VPWR VPWR _13196_/A sky130_fd_sc_hd__buf_1
XFILLER_120_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13968_ _13968_/A _13967_/X VGND VGND VPWR VPWR _13968_/X sky130_fd_sc_hd__or2b_1
XFILLER_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15707_ _15552_/A _14928_/B _14928_/Y VGND VGND VPWR VPWR _15707_/X sky130_fd_sc_hd__o21a_1
X_12919_ _12836_/X _12916_/Y _12917_/Y _12918_/X VGND VGND VPWR VPWR _12922_/B sky130_fd_sc_hd__o22a_1
XFILLER_19_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13899_ _13854_/X _13898_/Y _13854_/X _13898_/Y VGND VGND VPWR VPWR _13955_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15638_ _15671_/A _15671_/B VGND VGND VPWR VPWR _15638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15569_ _15429_/X _15568_/X _15429_/X _15568_/X VGND VGND VPWR VPWR _15655_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09090_ _09701_/A VGND VGND VPWR VPWR _09421_/A sky130_fd_sc_hd__buf_1
XFILLER_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09992_ _09992_/A _09993_/B VGND VGND VPWR VPWR _09992_/Y sky130_fd_sc_hd__nor2_1
X_08943_ _08939_/Y _11407_/A _08942_/Y VGND VGND VPWR VPWR _08952_/A sky130_fd_sc_hd__o21ai_1
XFILLER_96_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08874_ _08873_/Y _08867_/X _08873_/Y _08867_/X VGND VGND VPWR VPWR _08984_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09426_ _09426_/A _09433_/B VGND VGND VPWR VPWR _09426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09357_ _08694_/A _09862_/A _09348_/Y _09356_/X VGND VGND VPWR VPWR _09357_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08308_ _08308_/A VGND VGND VPWR VPWR _08308_/Y sky130_fd_sc_hd__inv_2
X_09288_ _09237_/A _09287_/Y _09237_/A _09287_/Y VGND VGND VPWR VPWR _10402_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08239_ _08239_/A VGND VGND VPWR VPWR _08239_/Y sky130_fd_sc_hd__inv_4
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11250_ _14047_/A _11252_/B VGND VGND VPWR VPWR _11250_/X sky130_fd_sc_hd__and2_1
XFILLER_133_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10201_ _10213_/A _10213_/B VGND VGND VPWR VPWR _10201_/Y sky130_fd_sc_hd__nor2_1
X_11181_ _11181_/A VGND VGND VPWR VPWR _11181_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10132_ _10132_/A _10132_/B VGND VGND VPWR VPWR _10133_/B sky130_fd_sc_hd__or2_1
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14940_ _14841_/A _14841_/B _14838_/X _14841_/Y VGND VGND VPWR VPWR _14940_/X sky130_fd_sc_hd__o2bb2a_1
X_10063_ _10063_/A _10063_/B VGND VGND VPWR VPWR _10063_/X sky130_fd_sc_hd__or2_1
X_14871_ _15548_/A _14924_/B VGND VGND VPWR VPWR _14871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13822_ _13759_/X _13821_/X _13759_/X _13821_/X VGND VGND VPWR VPWR _13843_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13753_ _13753_/A _13753_/B VGND VGND VPWR VPWR _13754_/A sky130_fd_sc_hd__or2_1
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10965_ _10962_/Y _12691_/A _10813_/X _10964_/Y VGND VGND VPWR VPWR _10965_/X sky130_fd_sc_hd__o22a_1
X_12704_ _12704_/A _12704_/B VGND VGND VPWR VPWR _12704_/X sky130_fd_sc_hd__and2_1
XFILLER_16_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16472_ _16472_/D _16456_/LO VGND VGND VPWR VPWR _16472_/Q sky130_fd_sc_hd__dlxtn_1
X_13684_ _13683_/A _13683_/B _11961_/X _13683_/X VGND VGND VPWR VPWR _13685_/A sky130_fd_sc_hd__o22a_1
X_10896_ _10896_/A VGND VGND VPWR VPWR _10896_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12635_ _14183_/A _12633_/X _12634_/X VGND VGND VPWR VPWR _12635_/X sky130_fd_sc_hd__o21a_1
X_15423_ _15356_/Y _15421_/Y _15422_/Y VGND VGND VPWR VPWR _15423_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12566_ _12566_/A VGND VGND VPWR VPWR _12566_/Y sky130_fd_sc_hd__inv_2
X_15354_ _15293_/X _15352_/X _15357_/B VGND VGND VPWR VPWR _15354_/X sky130_fd_sc_hd__o21a_1
X_14305_ _15966_/A _14395_/B VGND VGND VPWR VPWR _14305_/X sky130_fd_sc_hd__and2_1
X_11517_ _12376_/A VGND VGND VPWR VPWR _12685_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12497_ _12494_/Y _12495_/Y _12496_/Y VGND VGND VPWR VPWR _12497_/X sky130_fd_sc_hd__o21a_1
X_15285_ _15285_/A _15285_/B VGND VGND VPWR VPWR _15287_/B sky130_fd_sc_hd__and2_1
X_14236_ _14236_/A VGND VGND VPWR VPWR _14242_/A sky130_fd_sc_hd__inv_2
X_11448_ _12346_/A VGND VGND VPWR VPWR _15534_/A sky130_fd_sc_hd__buf_1
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14167_ _13447_/A _14144_/A _14142_/Y VGND VGND VPWR VPWR _14167_/Y sky130_fd_sc_hd__a21oi_1
X_11379_ _12311_/A _11379_/B VGND VGND VPWR VPWR _11379_/Y sky130_fd_sc_hd__nand2_1
X_13118_ _13062_/Y _13116_/X _13117_/Y VGND VGND VPWR VPWR _13118_/X sky130_fd_sc_hd__o21a_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _15461_/A _14031_/B _14031_/A _14031_/B VGND VGND VPWR VPWR _14098_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13774_/A VGND VGND VPWR VPWR _15240_/A sky130_fd_sc_hd__buf_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08590_ _09455_/B VGND VGND VPWR VPWR _09551_/A sky130_fd_sc_hd__buf_1
XFILLER_47_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09211_ _09553_/A _09731_/A VGND VGND VPWR VPWR _09212_/A sky130_fd_sc_hd__or2_1
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09142_ _09138_/Y _09140_/Y _09141_/Y VGND VGND VPWR VPWR _09175_/B sky130_fd_sc_hd__o21ai_1
X_09073_ _10016_/B _09073_/B VGND VGND VPWR VPWR _09074_/B sky130_fd_sc_hd__or2_1
XFILLER_131_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09975_ _09975_/A _09975_/B VGND VGND VPWR VPWR _09975_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08926_ _09817_/A VGND VGND VPWR VPWR _10102_/A sky130_fd_sc_hd__inv_2
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08857_ _10103_/A _08855_/Y _08916_/A _09460_/A VGND VGND VPWR VPWR _08857_/X sky130_fd_sc_hd__o22a_1
XFILLER_85_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08788_ _08712_/A _09470_/B _08712_/Y VGND VGND VPWR VPWR _08789_/A sky130_fd_sc_hd__a21oi_2
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10750_ _09952_/A _09631_/B _09632_/A VGND VGND VPWR VPWR _10751_/A sky130_fd_sc_hd__o21ai_1
XFILLER_111_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10681_ _10968_/A _10681_/B VGND VGND VPWR VPWR _10682_/A sky130_fd_sc_hd__or2_1
X_09409_ _09409_/A _09409_/B VGND VGND VPWR VPWR _09409_/Y sky130_fd_sc_hd__nor2_1
X_12420_ _12683_/A _12420_/B VGND VGND VPWR VPWR _12420_/X sky130_fd_sc_hd__or2_1
XFILLER_40_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12351_ _12351_/A _12351_/B VGND VGND VPWR VPWR _12351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11302_ _12946_/A VGND VGND VPWR VPWR _13780_/A sky130_fd_sc_hd__inv_2
X_15070_ _15070_/A _15036_/X VGND VGND VPWR VPWR _15070_/X sky130_fd_sc_hd__or2b_1
X_12282_ _12262_/X _12281_/X _12262_/X _12281_/X VGND VGND VPWR VPWR _12367_/B sky130_fd_sc_hd__a2bb2o_1
X_11233_ _14809_/A VGND VGND VPWR VPWR _12229_/A sky130_fd_sc_hd__inv_2
X_14021_ _15408_/A _13949_/B _13949_/Y VGND VGND VPWR VPWR _14021_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11164_ _12189_/A _11297_/B VGND VGND VPWR VPWR _11164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15972_ _15972_/A _15972_/B VGND VGND VPWR VPWR _15993_/B sky130_fd_sc_hd__or2_1
XFILLER_95_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11095_ _11186_/A _11093_/X _11094_/X VGND VGND VPWR VPWR _11095_/X sky130_fd_sc_hd__o21a_1
X_10115_ _10115_/A _10115_/B VGND VGND VPWR VPWR _10116_/A sky130_fd_sc_hd__or2_1
XFILLER_121_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14923_ _14875_/Y _14921_/X _14922_/Y VGND VGND VPWR VPWR _14923_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10046_ _10046_/A _10081_/B VGND VGND VPWR VPWR _10046_/X sky130_fd_sc_hd__and2_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14854_ _15353_/A _14958_/B VGND VGND VPWR VPWR _14854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14785_ _14735_/X _14784_/X _14735_/X _14784_/X VGND VGND VPWR VPWR _14786_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13805_ _14409_/A _13855_/B VGND VGND VPWR VPWR _13805_/Y sky130_fd_sc_hd__nor2_1
X_11997_ _10826_/A _11996_/A _10826_/Y _12084_/B VGND VGND VPWR VPWR _11999_/B sky130_fd_sc_hd__o22a_1
X_13736_ _13693_/X _13735_/X _13693_/X _13735_/X VGND VGND VPWR VPWR _13764_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10948_ _10948_/A VGND VGND VPWR VPWR _10948_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16455_ _16471_/Q _08230_/A _08233_/A _16392_/C _16343_/A VGND VGND VPWR VPWR _16471_/D
+ sky130_fd_sc_hd__o221a_2
X_15406_ _15406_/A _15406_/B VGND VGND VPWR VPWR _15406_/X sky130_fd_sc_hd__or2_1
X_13667_ _15134_/A _13625_/B _13625_/Y VGND VGND VPWR VPWR _13667_/Y sky130_fd_sc_hd__o21ai_1
X_10879_ _10879_/A _09412_/X VGND VGND VPWR VPWR _10880_/A sky130_fd_sc_hd__or2b_1
XFILLER_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16386_ _16058_/X _16386_/B VGND VGND VPWR VPWR _16386_/X sky130_fd_sc_hd__and2b_1
X_12618_ _12618_/A _12618_/B VGND VGND VPWR VPWR _12618_/X sky130_fd_sc_hd__or2_1
X_13598_ _13624_/A _13625_/B VGND VGND VPWR VPWR _13598_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12549_ _12549_/A VGND VGND VPWR VPWR _12549_/Y sky130_fd_sc_hd__inv_2
X_15337_ _15337_/A _15337_/B VGND VGND VPWR VPWR _15337_/X sky130_fd_sc_hd__or2_1
XFILLER_129_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15268_ _15268_/A _15216_/X VGND VGND VPWR VPWR _15268_/X sky130_fd_sc_hd__or2b_1
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 _08299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14219_ _14219_/A _12622_/X VGND VGND VPWR VPWR _14219_/X sky130_fd_sc_hd__or2b_1
XFILLER_125_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15199_ _15199_/A _15199_/B VGND VGND VPWR VPWR _15199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _09760_/A VGND VGND VPWR VPWR _09782_/A sky130_fd_sc_hd__inv_2
XFILLER_100_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08711_ _08711_/A _09472_/B VGND VGND VPWR VPWR _08711_/Y sky130_fd_sc_hd__nor2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _08618_/X _09693_/B _08618_/X _09693_/B VGND VGND VPWR VPWR _09692_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08642_ _08642_/A VGND VGND VPWR VPWR _08718_/A sky130_fd_sc_hd__inv_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer24 _14258_/A VGND VGND VPWR VPWR _14337_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer46 _09749_/X VGND VGND VPWR VPWR _11605_/A1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer35 _10190_/X VGND VGND VPWR VPWR _11325_/A1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer13 rebuffer14/X VGND VGND VPWR VPWR rebuffer13/X sky130_fd_sc_hd__dlygate4sd1_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08573_ _08573_/A VGND VGND VPWR VPWR _08573_/Y sky130_fd_sc_hd__inv_2
Xrebuffer57 _08398_/A VGND VGND VPWR VPWR rebuffer57/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09125_ _09421_/A _09126_/B VGND VGND VPWR VPWR _09125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09056_ _08781_/Y _09052_/A _08781_/A _09052_/Y VGND VGND VPWR VPWR _10012_/B sky130_fd_sc_hd__o22a_1
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09958_ _09958_/A _09958_/B VGND VGND VPWR VPWR _09958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08909_ _08683_/X _08908_/X _08683_/X _08908_/X VGND VGND VPWR VPWR _08970_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09889_ _09874_/X _09888_/X _09874_/X _09888_/X VGND VGND VPWR VPWR _09932_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11920_ _11987_/A VGND VGND VPWR VPWR _12776_/A sky130_fd_sc_hd__buf_1
XFILLER_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11851_ _11851_/A VGND VGND VPWR VPWR _11851_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14570_ _15270_/A _14571_/B VGND VGND VPWR VPWR _14570_/Y sky130_fd_sc_hd__nor2_1
X_11782_ _11731_/B _11781_/Y _11731_/B _11781_/Y VGND VGND VPWR VPWR _11783_/B sky130_fd_sc_hd__o2bb2a_1
X_10802_ _10801_/A _10801_/B _10801_/Y _09392_/A VGND VGND VPWR VPWR _10953_/A sky130_fd_sc_hd__o211a_1
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10733_ _11972_/A _10733_/B VGND VGND VPWR VPWR _10733_/Y sky130_fd_sc_hd__nand2_1
X_13521_ _13521_/A _13521_/B VGND VGND VPWR VPWR _13521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16240_ _16249_/A _16316_/A VGND VGND VPWR VPWR _16240_/Y sky130_fd_sc_hd__nor2_1
X_13452_ _13451_/Y _13307_/X _13209_/Y VGND VGND VPWR VPWR _13452_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10664_ _10664_/A _10664_/B VGND VGND VPWR VPWR _10664_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16171_ _16073_/X _16171_/B VGND VGND VPWR VPWR _16171_/X sky130_fd_sc_hd__and2b_1
X_13383_ _14131_/A _13443_/B VGND VGND VPWR VPWR _13383_/Y sky130_fd_sc_hd__nor2_1
X_12403_ _13544_/A _12404_/B VGND VGND VPWR VPWR _12403_/X sky130_fd_sc_hd__and2_1
X_10595_ _10530_/X _10594_/Y _10530_/X _10594_/Y VGND VGND VPWR VPWR _10642_/B sky130_fd_sc_hd__a2bb2o_1
X_12334_ _14032_/A _12226_/B _12226_/Y VGND VGND VPWR VPWR _12334_/Y sky130_fd_sc_hd__o21ai_1
X_15122_ _15122_/A _15122_/B VGND VGND VPWR VPWR _15122_/Y sky130_fd_sc_hd__nand2_1
X_15053_ _15047_/X _15052_/Y _15047_/X _15052_/Y VGND VGND VPWR VPWR _15054_/B sky130_fd_sc_hd__a2bb2o_1
X_14004_ _13960_/X _14003_/Y _13960_/X _14003_/Y VGND VGND VPWR VPWR _14065_/B sky130_fd_sc_hd__a2bb2o_1
X_12265_ _12263_/A _12263_/B _12263_/X _12264_/Y VGND VGND VPWR VPWR _12371_/B sky130_fd_sc_hd__a22o_1
XFILLER_5_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11216_ _12220_/A VGND VGND VPWR VPWR _14027_/A sky130_fd_sc_hd__buf_1
X_12196_ _12195_/A _12254_/B _12195_/Y VGND VGND VPWR VPWR _12196_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11147_ _11147_/A VGND VGND VPWR VPWR _11147_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15955_ _15936_/X _15953_/X _16014_/B VGND VGND VPWR VPWR _15955_/X sky130_fd_sc_hd__o21a_1
X_11078_ _15392_/A _11078_/B VGND VGND VPWR VPWR _11078_/X sky130_fd_sc_hd__or2_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15886_ _15886_/A _15886_/B VGND VGND VPWR VPWR _15886_/Y sky130_fd_sc_hd__nand2_1
X_14906_ _14906_/A _14906_/B VGND VGND VPWR VPWR _14906_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10029_ _09331_/A _09331_/B _10038_/B _10028_/X VGND VGND VPWR VPWR _10029_/X sky130_fd_sc_hd__o22a_1
XFILLER_91_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14837_ _14757_/A _14757_/B _14750_/X _14757_/Y VGND VGND VPWR VPWR _14837_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14768_ _15351_/A _14830_/B _14767_/Y VGND VGND VPWR VPWR _14768_/Y sky130_fd_sc_hd__o21ai_1
X_14699_ _15341_/A _14655_/B _14655_/Y VGND VGND VPWR VPWR _14699_/Y sky130_fd_sc_hd__o21ai_1
X_13719_ _13719_/A _13719_/B VGND VGND VPWR VPWR _13720_/B sky130_fd_sc_hd__or2_1
X_16438_ _16460_/Q _16459_/Q _16458_/Q _16447_/B _16437_/X VGND VGND VPWR VPWR _16438_/X
+ sky130_fd_sc_hd__o41a_1
X_16369_ _16324_/A _16324_/B _16324_/Y VGND VGND VPWR VPWR _16369_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09812_ _08819_/A _08610_/A _09456_/Y _09811_/X VGND VGND VPWR VPWR _09812_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09743_ _09743_/A _09743_/B VGND VGND VPWR VPWR _09743_/X sky130_fd_sc_hd__or2_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09674_ _09655_/X _09673_/X _09655_/X _09673_/X VGND VGND VPWR VPWR _09675_/B sky130_fd_sc_hd__a2bb2oi_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08625_ _08625_/A VGND VGND VPWR VPWR _08625_/Y sky130_fd_sc_hd__clkinvlp_2
Xclkbuf_1_0__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _08229_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_82_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08556_ _09859_/A VGND VGND VPWR VPWR _09737_/A sky130_fd_sc_hd__inv_2
XFILLER_23_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08487_ _08266_/A _08346_/B _08477_/Y _08599_/A VGND VGND VPWR VPWR _08587_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09108_ _09539_/B _09030_/B _09031_/B VGND VGND VPWR VPWR _09108_/Y sky130_fd_sc_hd__a21boi_1
X_10380_ _11808_/A _10452_/B _10379_/Y VGND VGND VPWR VPWR _10381_/A sky130_fd_sc_hd__o21ai_2
XFILLER_124_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09039_ _09529_/B _09038_/B _09155_/B VGND VGND VPWR VPWR _09040_/A sky130_fd_sc_hd__a21bo_1
XFILLER_123_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12050_ _12045_/Y _12048_/Y _12049_/Y VGND VGND VPWR VPWR _12050_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11001_ _12103_/A _11000_/B _11000_/Y VGND VGND VPWR VPWR _11001_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_132_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15740_ _15752_/A _15740_/B VGND VGND VPWR VPWR _16110_/A sky130_fd_sc_hd__nor2_1
X_12952_ _14948_/A _12953_/B VGND VGND VPWR VPWR _12954_/A sky130_fd_sc_hd__and2_1
XFILLER_46_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15671_ _15671_/A _15671_/B VGND VGND VPWR VPWR _15671_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11903_ _11903_/A VGND VGND VPWR VPWR _11903_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14622_ _14622_/A VGND VGND VPWR VPWR _15339_/A sky130_fd_sc_hd__buf_1
XFILLER_61_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12883_ _12852_/X _12882_/Y _12852_/X _12882_/Y VGND VGND VPWR VPWR _12940_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _11794_/A _11794_/B _11794_/A _11794_/B VGND VGND VPWR VPWR _11834_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14553_ _14514_/X _14552_/X _14514_/X _14552_/X VGND VGND VPWR VPWR _14579_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11765_ _10381_/A _11764_/A _10381_/Y _11808_/B VGND VGND VPWR VPWR _11767_/B sky130_fd_sc_hd__o22a_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _12789_/A VGND VGND VPWR VPWR _13994_/A sky130_fd_sc_hd__buf_6
X_10716_ _13068_/A _10716_/B VGND VGND VPWR VPWR _10716_/Y sky130_fd_sc_hd__nand2_1
X_14484_ _14484_/A VGND VGND VPWR VPWR _15199_/A sky130_fd_sc_hd__buf_1
X_13504_ _13506_/A VGND VGND VPWR VPWR _15044_/A sky130_fd_sc_hd__buf_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16223_ _16223_/A VGND VGND VPWR VPWR _16223_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13435_ _14111_/A _13435_/B VGND VGND VPWR VPWR _13435_/Y sky130_fd_sc_hd__nand2_1
X_10647_ _10647_/A VGND VGND VPWR VPWR _10647_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer4 rebuffer5/X VGND VGND VPWR VPWR rebuffer4/X sky130_fd_sc_hd__dlygate4sd1_1
X_16154_ _16270_/A _16336_/A VGND VGND VPWR VPWR _16154_/Y sky130_fd_sc_hd__nor2_1
X_13366_ _13366_/A _13366_/B VGND VGND VPWR VPWR _13366_/X sky130_fd_sc_hd__or2_1
X_10578_ _10547_/X _10577_/X _10547_/X _10577_/X VGND VGND VPWR VPWR _10661_/B sky130_fd_sc_hd__a2bb2o_1
X_16085_ _16082_/Y _16233_/A _16084_/Y VGND VGND VPWR VPWR _16089_/B sky130_fd_sc_hd__o21ai_1
XFILLER_127_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12317_ _13404_/A VGND VGND VPWR VPWR _14081_/A sky130_fd_sc_hd__inv_2
X_13297_ _14738_/A _13297_/B VGND VGND VPWR VPWR _13297_/Y sky130_fd_sc_hd__nand2_1
X_15105_ _15103_/X _15105_/B VGND VGND VPWR VPWR _15105_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12248_ _14059_/A _12208_/B _12208_/Y _12247_/X VGND VGND VPWR VPWR _12248_/X sky130_fd_sc_hd__a2bb2o_1
X_15036_ _15036_/A _15036_/B VGND VGND VPWR VPWR _15036_/X sky130_fd_sc_hd__or2_1
XFILLER_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12179_ _11152_/A _12178_/A _11152_/Y _12270_/B VGND VGND VPWR VPWR _12181_/B sky130_fd_sc_hd__o22a_1
XFILLER_110_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15938_ _15889_/X _15937_/Y _15889_/X _15937_/Y VGND VGND VPWR VPWR _15952_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15869_ _15869_/A VGND VGND VPWR VPWR _15894_/A sky130_fd_sc_hd__inv_2
XFILLER_91_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08410_ _08409_/A _08354_/Y _08409_/Y _08354_/A _08419_/A VGND VGND VPWR VPWR _09225_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09390_ _10420_/B VGND VGND VPWR VPWR _09391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08341_ input30/X _08341_/B VGND VGND VPWR VPWR _08342_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08272_ _08272_/A input11/X VGND VGND VPWR VPWR _08364_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09726_ _09770_/A _09770_/B _09725_/Y VGND VGND VPWR VPWR _09727_/A sky130_fd_sc_hd__o21ai_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09657_ _09603_/Y _09655_/X _09656_/Y VGND VGND VPWR VPWR _09657_/X sky130_fd_sc_hd__o21a_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08716_/B VGND VGND VPWR VPWR _08610_/A sky130_fd_sc_hd__buf_1
X_09588_ _09989_/A VGND VGND VPWR VPWR _09990_/A sky130_fd_sc_hd__buf_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08539_ _08538_/A _08323_/Y _08538_/Y _08323_/A VGND VGND VPWR VPWR _08540_/B sky130_fd_sc_hd__o22a_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11550_ _12955_/A _11646_/B _11549_/Y VGND VGND VPWR VPWR _11550_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10501_ _12928_/A VGND VGND VPWR VPWR _11840_/A sky130_fd_sc_hd__inv_2
XFILLER_7_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13220_ _14771_/A _13303_/B VGND VGND VPWR VPWR _13220_/Y sky130_fd_sc_hd__nor2_1
X_11481_ _11482_/A VGND VGND VPWR VPWR _14744_/A sky130_fd_sc_hd__buf_1
XFILLER_7_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10432_ _10511_/A _10430_/X _10431_/X VGND VGND VPWR VPWR _10432_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13151_ _15243_/A _13119_/B _13119_/Y VGND VGND VPWR VPWR _13151_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10363_ _09971_/A _10362_/Y _09971_/Y _10362_/A _10445_/A VGND VGND VPWR VPWR _11758_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13082_ _15258_/A _13109_/B VGND VGND VPWR VPWR _13082_/Y sky130_fd_sc_hd__nor2_1
X_12102_ _12163_/A _12101_/Y _12163_/A _12101_/Y VGND VGND VPWR VPWR _12160_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12033_ _12055_/A VGND VGND VPWR VPWR _13188_/A sky130_fd_sc_hd__buf_1
X_10294_ _10335_/B VGND VGND VPWR VPWR _10294_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15723_ _15685_/A _15685_/B _15685_/Y VGND VGND VPWR VPWR _15723_/Y sky130_fd_sc_hd__o21ai_1
X_13984_ _13984_/A _13984_/B VGND VGND VPWR VPWR _13985_/B sky130_fd_sc_hd__or2_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12935_ _12896_/Y _12933_/X _12934_/Y VGND VGND VPWR VPWR _12935_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15654_ _15667_/A _15667_/B VGND VGND VPWR VPWR _15654_/X sky130_fd_sc_hd__and2_1
X_12866_ _13872_/A _12861_/B _12861_/Y VGND VGND VPWR VPWR _12866_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15585_ _15685_/A _15685_/B VGND VGND VPWR VPWR _15585_/Y sky130_fd_sc_hd__nor2_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14590_/X _14604_/X _14590_/X _14604_/X VGND VGND VPWR VPWR _14664_/B sky130_fd_sc_hd__a2bb2o_1
X_11817_ _12772_/A _11851_/A _11816_/Y VGND VGND VPWR VPWR _11817_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _14536_/A _14535_/X VGND VGND VPWR VPWR _14536_/X sky130_fd_sc_hd__or2b_1
X_12797_ _12782_/A _12782_/B _12782_/Y VGND VGND VPWR VPWR _12797_/Y sky130_fd_sc_hd__o21ai_1
X_11748_ _11748_/A _11748_/B VGND VGND VPWR VPWR _11748_/X sky130_fd_sc_hd__or2_1
XFILLER_14_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14467_ _14444_/Y _14465_/X _14466_/Y VGND VGND VPWR VPWR _14467_/X sky130_fd_sc_hd__o21a_1
X_11679_ _11620_/Y _11624_/Y _12428_/A _11618_/A VGND VGND VPWR VPWR _11679_/X sky130_fd_sc_hd__a2bb2o_2
X_16206_ _16104_/A _15805_/B _15805_/Y VGND VGND VPWR VPWR _16208_/A sky130_fd_sc_hd__o21ai_1
X_14398_ _14282_/X _14398_/B VGND VGND VPWR VPWR _14398_/Y sky130_fd_sc_hd__nand2b_1
X_13418_ _13340_/A _13340_/B _13340_/A _13340_/B VGND VGND VPWR VPWR _13418_/X sky130_fd_sc_hd__a2bb2o_1
X_16137_ _16136_/A _16136_/B _16136_/X VGND VGND VPWR VPWR _16137_/Y sky130_fd_sc_hd__a21boi_1
X_13349_ _13349_/A VGND VGND VPWR VPWR _13349_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16068_ _16044_/A _16044_/B _16044_/Y VGND VGND VPWR VPWR _16068_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15019_ _11768_/Y _15000_/X _11768_/Y _15000_/X VGND VGND VPWR VPWR _15034_/B sky130_fd_sc_hd__a2bb2o_1
X_08890_ _08978_/A _08978_/B VGND VGND VPWR VPWR _08890_/X sky130_fd_sc_hd__and2_1
XFILLER_111_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09511_ _09494_/A _09494_/B _09494_/Y _09510_/X VGND VGND VPWR VPWR _09511_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09442_ _09198_/X _09359_/X _09198_/X _09359_/X VGND VGND VPWR VPWR _09442_/X sky130_fd_sc_hd__o2bb2a_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09373_ _09373_/A VGND VGND VPWR VPWR _09431_/B sky130_fd_sc_hd__inv_2
XFILLER_40_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08324_ _08324_/A VGND VGND VPWR VPWR _08324_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08255_ input16/X VGND VGND VPWR VPWR _08331_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10981_ _10967_/X _10980_/Y _10967_/X _10980_/Y VGND VGND VPWR VPWR _11138_/A sky130_fd_sc_hd__o2bb2a_1
X_09709_ _09709_/A _09709_/B VGND VGND VPWR VPWR _09709_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12720_ _12685_/A _12685_/B _12685_/Y _12719_/X VGND VGND VPWR VPWR _12720_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12651_ _12651_/A _12651_/B VGND VGND VPWR VPWR _14162_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11602_ _11602_/A _11602_/B VGND VGND VPWR VPWR _11602_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12582_ _14910_/A _12336_/B _12336_/Y VGND VGND VPWR VPWR _12583_/A sky130_fd_sc_hd__o21ai_1
X_15370_ _15344_/X _15369_/X _15344_/X _15369_/X VGND VGND VPWR VPWR _15412_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14321_ _15863_/A _14268_/B _14268_/Y VGND VGND VPWR VPWR _14321_/Y sky130_fd_sc_hd__o21ai_1
X_11533_ _11533_/A VGND VGND VPWR VPWR _11533_/Y sky130_fd_sc_hd__clkinvlp_2
X_14252_ _14252_/A VGND VGND VPWR VPWR _14252_/Y sky130_fd_sc_hd__inv_2
X_11464_ _11572_/A _11464_/B VGND VGND VPWR VPWR _12410_/A sky130_fd_sc_hd__or2_2
XFILLER_99_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13203_ _13150_/Y _13201_/X _13202_/Y VGND VGND VPWR VPWR _13203_/X sky130_fd_sc_hd__o21a_1
X_10415_ _12826_/A _10431_/B VGND VGND VPWR VPWR _10511_/A sky130_fd_sc_hd__and2_1
XFILLER_109_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14183_ _14183_/A _12634_/X VGND VGND VPWR VPWR _14183_/X sky130_fd_sc_hd__or2b_1
X_11395_ _11395_/A VGND VGND VPWR VPWR _11395_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13134_ _13966_/A VGND VGND VPWR VPWR _15167_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10346_ _10906_/A _10346_/B VGND VGND VPWR VPWR _10347_/A sky130_fd_sc_hd__or2_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13065_ _13065_/A _13025_/X VGND VGND VPWR VPWR _13065_/X sky130_fd_sc_hd__or2b_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ _10277_/A VGND VGND VPWR VPWR _10277_/Y sky130_fd_sc_hd__inv_2
X_12016_ _13198_/A _12065_/B VGND VGND VPWR VPWR _12016_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13967_ _15167_/A _13967_/B VGND VGND VPWR VPWR _13967_/X sky130_fd_sc_hd__or2_1
XFILLER_19_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15706_ _16125_/A _15823_/B VGND VGND VPWR VPWR _15706_/X sky130_fd_sc_hd__and2_1
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12918_ _12837_/A _12837_/B _12837_/X VGND VGND VPWR VPWR _12918_/X sky130_fd_sc_hd__o21ba_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15637_ _14380_/X _15636_/Y _14380_/X _15636_/Y VGND VGND VPWR VPWR _15671_/B sky130_fd_sc_hd__a2bb2o_1
X_13898_ _14409_/A _13855_/B _13855_/Y VGND VGND VPWR VPWR _13898_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12849_ _12849_/A _12849_/B VGND VGND VPWR VPWR _12849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _15562_/X _15567_/Y _15562_/X _15567_/Y VGND VGND VPWR VPWR _15568_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15499_ _15482_/X _15498_/X _15482_/X _15498_/X VGND VGND VPWR VPWR _15546_/B sky130_fd_sc_hd__a2bb2o_1
X_14519_ _15196_/A _14519_/B VGND VGND VPWR VPWR _14519_/X sky130_fd_sc_hd__or2_1
XFILLER_115_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09991_ _09967_/Y _09989_/Y _09990_/Y VGND VGND VPWR VPWR _09993_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08942_ _08942_/A _08942_/B VGND VGND VPWR VPWR _08942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08873_ _08762_/A _10133_/A _08762_/Y VGND VGND VPWR VPWR _08873_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09425_ _09265_/A _09423_/Y _09424_/Y VGND VGND VPWR VPWR _09433_/B sky130_fd_sc_hd__o21ai_1
XFILLER_40_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09356_ _08692_/A _09861_/A _09350_/Y _09355_/X VGND VGND VPWR VPWR _09356_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08307_ _08307_/A _08307_/B VGND VGND VPWR VPWR _08308_/A sky130_fd_sc_hd__or2_1
X_09287_ _09230_/A _09800_/A _09230_/Y VGND VGND VPWR VPWR _09287_/Y sky130_fd_sc_hd__a21oi_1
X_08238_ _08238_/A _08238_/B VGND VGND VPWR VPWR _08239_/A sky130_fd_sc_hd__or2_2
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10200_ _10108_/A _10109_/A _10108_/Y _10109_/Y _10346_/B VGND VGND VPWR VPWR _10213_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11180_ _09436_/A _09141_/B _09141_/Y VGND VGND VPWR VPWR _11181_/A sky130_fd_sc_hd__o21ai_1
XFILLER_133_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10131_ _10131_/A _10131_/B VGND VGND VPWR VPWR _10132_/B sky130_fd_sc_hd__or2_1
XFILLER_121_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10062_ _10020_/X _10061_/Y _10020_/X _10061_/Y VGND VGND VPWR VPWR _10063_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14870_ _14825_/X _14869_/X _14825_/X _14869_/X VGND VGND VPWR VPWR _14924_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13821_ _13821_/A _13760_/X VGND VGND VPWR VPWR _13821_/X sky130_fd_sc_hd__or2b_1
XFILLER_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13752_ _13752_/A _13752_/B VGND VGND VPWR VPWR _13752_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12703_ _10226_/X _12658_/Y _10226_/X _12658_/Y VGND VGND VPWR VPWR _12704_/B sky130_fd_sc_hd__a2bb2o_1
X_10964_ _10964_/A _11999_/A VGND VGND VPWR VPWR _10964_/Y sky130_fd_sc_hd__nor2_1
X_16471_ _08229_/A _16471_/D VGND VGND VPWR VPWR _16471_/Q sky130_fd_sc_hd__dfxtp_1
X_13683_ _13683_/A _13683_/B VGND VGND VPWR VPWR _13683_/X sky130_fd_sc_hd__and2_1
XFILLER_16_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10895_ _10895_/A _09407_/X VGND VGND VPWR VPWR _10896_/A sky130_fd_sc_hd__or2b_1
X_12634_ _12634_/A _12634_/B VGND VGND VPWR VPWR _12634_/X sky130_fd_sc_hd__or2_1
X_15422_ _15422_/A _15422_/B VGND VGND VPWR VPWR _15422_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12565_ _12626_/A _12626_/B VGND VGND VPWR VPWR _14207_/A sky130_fd_sc_hd__and2_1
X_15353_ _15353_/A _15353_/B VGND VGND VPWR VPWR _15357_/B sky130_fd_sc_hd__or2_1
XFILLER_8_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14304_ _14275_/Y _14303_/Y _14275_/Y _14303_/Y VGND VGND VPWR VPWR _14395_/B sky130_fd_sc_hd__a2bb2o_1
X_11516_ _11519_/A VGND VGND VPWR VPWR _11516_/Y sky130_fd_sc_hd__inv_2
X_12496_ _12496_/A _12496_/B VGND VGND VPWR VPWR _12496_/Y sky130_fd_sc_hd__nand2_1
X_15284_ _14953_/A _15234_/B _15234_/Y _15283_/X VGND VGND VPWR VPWR _15284_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_11_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14235_ _14235_/A _15839_/A VGND VGND VPWR VPWR _14236_/A sky130_fd_sc_hd__or2_1
X_11447_ _11257_/X _11446_/Y _11257_/X _11446_/Y VGND VGND VPWR VPWR _12556_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14166_ _14164_/X _14166_/B VGND VGND VPWR VPWR _14166_/Y sky130_fd_sc_hd__nand2b_1
X_11378_ _11260_/X _11377_/Y _11260_/X _11377_/Y VGND VGND VPWR VPWR _11379_/B sky130_fd_sc_hd__a2bb2o_1
X_13117_ _15246_/A _13117_/B VGND VGND VPWR VPWR _13117_/Y sky130_fd_sc_hd__nand2_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _09955_/A _09955_/B _09955_/X VGND VGND VPWR VPWR _10330_/A sky130_fd_sc_hd__o21ba_1
XFILLER_112_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14097_ _14097_/A _14100_/B VGND VGND VPWR VPWR _14097_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13048_/A VGND VGND VPWR VPWR _13774_/A sky130_fd_sc_hd__inv_2
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14999_ _12704_/A _11746_/Y _11739_/Y _14998_/X VGND VGND VPWR VPWR _14999_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09210_ _09857_/A VGND VGND VPWR VPWR _09731_/A sky130_fd_sc_hd__inv_2
X_09141_ _09436_/A _09141_/B VGND VGND VPWR VPWR _09141_/Y sky130_fd_sc_hd__nand2_1
X_09072_ _10017_/B _09072_/B VGND VGND VPWR VPWR _09073_/B sky130_fd_sc_hd__or2_1
XFILLER_128_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09974_ _09974_/A _09975_/B VGND VGND VPWR VPWR _09974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08925_ _08930_/A _09541_/A VGND VGND VPWR VPWR _09817_/A sky130_fd_sc_hd__or2_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08856_ _08856_/A _08856_/B VGND VGND VPWR VPWR _09460_/A sky130_fd_sc_hd__or2_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08787_ _09323_/A VGND VGND VPWR VPWR _09490_/A sky130_fd_sc_hd__buf_1
XFILLER_25_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10680_ _10076_/X _10679_/X _10076_/X _10679_/X VGND VGND VPWR VPWR _10681_/B sky130_fd_sc_hd__a2bb2o_1
X_09408_ _09296_/A _10895_/A _09407_/X VGND VGND VPWR VPWR _09409_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09339_ _08753_/Y _09337_/Y _09338_/X VGND VGND VPWR VPWR _09339_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12350_ _12244_/X _12349_/Y _12244_/X _12349_/Y VGND VGND VPWR VPWR _12551_/A sky130_fd_sc_hd__a2bb2o_1
X_12281_ _11275_/A _12369_/B _11275_/A _12369_/B VGND VGND VPWR VPWR _12281_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11301_ _11299_/Y _11300_/Y _11300_/B _09927_/B _10794_/X VGND VGND VPWR VPWR _12946_/A
+ sky130_fd_sc_hd__o221a_2
X_11232_ _11232_/A _11251_/B VGND VGND VPWR VPWR _14809_/A sky130_fd_sc_hd__or2_1
X_14020_ _14020_/A _14055_/B VGND VGND VPWR VPWR _14076_/A sky130_fd_sc_hd__and2_1
XFILLER_122_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11163_ _11129_/X _11162_/X _11129_/X _11162_/X VGND VGND VPWR VPWR _11297_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10114_ _10114_/A _10114_/B VGND VGND VPWR VPWR _10115_/A sky130_fd_sc_hd__or2_1
X_15971_ _15918_/Y _15969_/Y _15970_/Y VGND VGND VPWR VPWR _15971_/X sky130_fd_sc_hd__o21a_1
X_11094_ _13897_/A _11094_/B VGND VGND VPWR VPWR _11094_/X sky130_fd_sc_hd__or2_1
XFILLER_76_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14922_ _15546_/A _14922_/B VGND VGND VPWR VPWR _14922_/Y sky130_fd_sc_hd__nand2_1
X_10045_ _10026_/X _10044_/Y _10026_/X _10044_/Y VGND VGND VPWR VPWR _10081_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14853_ _14834_/X _14852_/Y _14834_/X _14852_/Y VGND VGND VPWR VPWR _14958_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13804_ _13771_/X _13803_/X _13771_/X _13803_/X VGND VGND VPWR VPWR _13855_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14784_ _14784_/A _14736_/X VGND VGND VPWR VPWR _14784_/X sky130_fd_sc_hd__or2b_1
X_11996_ _11996_/A VGND VGND VPWR VPWR _12084_/B sky130_fd_sc_hd__inv_2
X_13735_ _13735_/A _13694_/X VGND VGND VPWR VPWR _13735_/X sky130_fd_sc_hd__or2b_1
X_10947_ _10946_/Y _10792_/X _10839_/Y VGND VGND VPWR VPWR _10947_/X sky130_fd_sc_hd__o21a_1
X_16454_ _16454_/A _16454_/B _16404_/B VGND VGND VPWR VPWR _16454_/Y sky130_fd_sc_hd__nor3b_1
X_13666_ _13694_/A _13694_/B VGND VGND VPWR VPWR _13735_/A sky130_fd_sc_hd__and2_1
XFILLER_31_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12617_ _12617_/A VGND VGND VPWR VPWR _14235_/A sky130_fd_sc_hd__inv_2
X_15405_ _15459_/A _15403_/X _15404_/X VGND VGND VPWR VPWR _15405_/X sky130_fd_sc_hd__o21a_1
X_10878_ _10878_/A _10878_/B VGND VGND VPWR VPWR _10878_/X sky130_fd_sc_hd__and2_1
XFILLER_129_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16385_ _16136_/A _16136_/B _16136_/X _16274_/Y VGND VGND VPWR VPWR _16385_/X sky130_fd_sc_hd__a22o_1
X_13597_ _13576_/X _13596_/Y _13576_/X _13596_/Y VGND VGND VPWR VPWR _13625_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12548_ _14916_/A _11455_/B _11455_/Y VGND VGND VPWR VPWR _12549_/A sky130_fd_sc_hd__o21ai_1
X_15336_ _15384_/A _15334_/X _15335_/X VGND VGND VPWR VPWR _15336_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12479_ _12403_/X _12359_/X _12405_/B VGND VGND VPWR VPWR _12479_/Y sky130_fd_sc_hd__o21ai_2
X_15267_ _15272_/A _15272_/B VGND VGND VPWR VPWR _15324_/A sky130_fd_sc_hd__and2_1
XANTENNA_2 _08299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14218_ _14230_/A _14218_/B VGND VGND VPWR VPWR _15875_/A sky130_fd_sc_hd__or2_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15198_ _15151_/X _15197_/Y _15151_/X _15197_/Y VGND VGND VPWR VPWR _15199_/B sky130_fd_sc_hd__a2bb2o_1
X_14149_ _14145_/X _14148_/Y _13449_/A _14148_/B VGND VGND VPWR VPWR _14149_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _08710_/A _09474_/B VGND VGND VPWR VPWR _08710_/Y sky130_fd_sc_hd__nor2_1
X_09690_ _09690_/A _09690_/B VGND VGND VPWR VPWR _09693_/B sky130_fd_sc_hd__or2_1
X_08641_ _08719_/B VGND VGND VPWR VPWR _09230_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer25 _08395_/A VGND VGND VPWR VPWR _08856_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer14 rebuffer15/X VGND VGND VPWR VPWR rebuffer14/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer36 _09748_/A VGND VGND VPWR VPWR _11599_/A1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer47 _12435_/Y VGND VGND VPWR VPWR _14973_/B1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer58 _11723_/B VGND VGND VPWR VPWR _11717_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_35_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08572_ _08572_/A _10116_/B VGND VGND VPWR VPWR _08573_/A sky130_fd_sc_hd__or2_1
XFILLER_35_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09124_ _09120_/Y _09122_/Y _09123_/Y VGND VGND VPWR VPWR _09126_/B sky130_fd_sc_hd__o21ai_1
X_09055_ _08773_/Y _09054_/A _08773_/A _09054_/Y VGND VGND VPWR VPWR _10011_/B sky130_fd_sc_hd__o22a_1
XFILLER_123_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09957_ _09957_/A _09958_/B VGND VGND VPWR VPWR _09957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08908_ _09549_/A _08609_/A _08611_/A VGND VGND VPWR VPWR _08908_/X sky130_fd_sc_hd__o21a_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09888_/A _09888_/B VGND VGND VPWR VPWR _09888_/X sky130_fd_sc_hd__or2_1
XFILLER_18_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08839_ _08839_/A VGND VGND VPWR VPWR _08839_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_18_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11850_ _11850_/A _11850_/B VGND VGND VPWR VPWR _11850_/X sky130_fd_sc_hd__or2_1
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11781_ _12766_/A _11780_/B _11780_/Y VGND VGND VPWR VPWR _11781_/Y sky130_fd_sc_hd__a21oi_1
X_10801_ _10801_/A _10801_/B VGND VGND VPWR VPWR _10801_/Y sky130_fd_sc_hd__nand2_1
X_10732_ _10641_/A _10731_/Y _10641_/A _10731_/Y VGND VGND VPWR VPWR _10733_/B sky130_fd_sc_hd__a2bb2o_1
X_13520_ _10388_/X _13483_/X _10388_/X _13483_/X VGND VGND VPWR VPWR _13521_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13451_ _14934_/A _13451_/B VGND VGND VPWR VPWR _13451_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10663_ _09268_/A _09268_/B _09268_/X VGND VGND VPWR VPWR _10664_/B sky130_fd_sc_hd__a21boi_1
XFILLER_13_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16170_ _16266_/A _16332_/A VGND VGND VPWR VPWR _16170_/Y sky130_fd_sc_hd__nor2_1
X_13382_ _13367_/X _13381_/X _13367_/X _13381_/X VGND VGND VPWR VPWR _13443_/B sky130_fd_sc_hd__a2bb2o_1
X_12402_ _12361_/X _12401_/Y _12361_/X _12401_/Y VGND VGND VPWR VPWR _12404_/B sky130_fd_sc_hd__a2bb2o_1
X_10594_ _13624_/A _10531_/B _10531_/Y VGND VGND VPWR VPWR _10594_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12333_ _13397_/A _12336_/B VGND VGND VPWR VPWR _12333_/Y sky130_fd_sc_hd__nor2_1
X_15121_ _15095_/X _15120_/Y _15095_/X _15120_/Y VGND VGND VPWR VPWR _15122_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15052_ _15050_/X _15052_/B VGND VGND VPWR VPWR _15052_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14003_ _15420_/A _13961_/B _13961_/Y VGND VGND VPWR VPWR _14003_/Y sky130_fd_sc_hd__o21ai_1
X_12264_ _12264_/A VGND VGND VPWR VPWR _12264_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11215_ _13334_/A VGND VGND VPWR VPWR _12220_/A sky130_fd_sc_hd__inv_2
X_12195_ _12195_/A _12254_/B VGND VGND VPWR VPWR _12195_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11146_ _10240_/B _10147_/B _10147_/Y VGND VGND VPWR VPWR _11147_/A sky130_fd_sc_hd__a21oi_1
X_15954_ _15954_/A _15954_/B VGND VGND VPWR VPWR _16014_/B sky130_fd_sc_hd__or2_1
X_11077_ _12139_/A VGND VGND VPWR VPWR _15392_/A sky130_fd_sc_hd__buf_1
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14905_ _14904_/A _14904_/B _12611_/A _14904_/Y VGND VGND VPWR VPWR _14905_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10028_ _09332_/A _09332_/B _10041_/B _10027_/X VGND VGND VPWR VPWR _10028_/X sky130_fd_sc_hd__o22a_1
X_15885_ _15885_/A _15885_/B VGND VGND VPWR VPWR _15885_/X sky130_fd_sc_hd__or2_1
XFILLER_91_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14836_ _14836_/A VGND VGND VPWR VPWR _15178_/A sky130_fd_sc_hd__buf_1
XFILLER_64_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14767_ _15351_/A _14830_/B VGND VGND VPWR VPWR _14767_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11979_ _11942_/Y _11977_/X _11978_/Y VGND VGND VPWR VPWR _11979_/X sky130_fd_sc_hd__o21a_1
X_13718_ _13719_/A _13719_/B VGND VGND VPWR VPWR _13718_/X sky130_fd_sc_hd__and2_1
XFILLER_44_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14698_ _14734_/A _14734_/B VGND VGND VPWR VPWR _14788_/A sky130_fd_sc_hd__and2_1
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16437_ _16467_/Q _16437_/B _16465_/Q _16437_/D VGND VGND VPWR VPWR _16437_/X sky130_fd_sc_hd__or4_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13649_ _13648_/A _13648_/B _13708_/A VGND VGND VPWR VPWR _13649_/Y sky130_fd_sc_hd__o21ai_1
X_16368_ _16357_/X _16463_/Q _16358_/X _16407_/A _16361_/X VGND VGND VPWR VPWR _16463_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_117_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15319_ _15274_/X _15318_/Y _15274_/X _15318_/Y VGND VGND VPWR VPWR _15335_/B sky130_fd_sc_hd__a2bb2o_1
X_16299_ _16326_/A _16326_/B VGND VGND VPWR VPWR _16299_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09811_ _08962_/X _08623_/A _09457_/Y _09810_/X VGND VGND VPWR VPWR _09811_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09742_ _09742_/A _09742_/B VGND VGND VPWR VPWR _09745_/A sky130_fd_sc_hd__or2_1
XFILLER_101_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09673_ _09984_/A _09656_/B _09656_/Y VGND VGND VPWR VPWR _09673_/X sky130_fd_sc_hd__o21a_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08624_ _08624_/A VGND VGND VPWR VPWR _08624_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08555_ _10011_/A _08555_/B VGND VGND VPWR VPWR _09859_/A sky130_fd_sc_hd__or2_2
XFILLER_70_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08486_ _08269_/A _08352_/B _08478_/Y _08612_/A VGND VGND VPWR VPWR _08599_/A sky130_fd_sc_hd__o22a_1
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09107_ _09714_/A _09107_/B VGND VGND VPWR VPWR _09107_/X sky130_fd_sc_hd__and2_1
XFILLER_109_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09038_ _09529_/B _09038_/B VGND VGND VPWR VPWR _09155_/B sky130_fd_sc_hd__or2_1
XFILLER_131_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11000_ _12103_/A _11000_/B VGND VGND VPWR VPWR _11000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12951_ _12865_/X _12950_/X _12865_/X _12950_/X VGND VGND VPWR VPWR _12953_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15670_ _15646_/Y _15668_/Y _15669_/Y VGND VGND VPWR VPWR _15670_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11902_ _11882_/Y _11900_/Y _11901_/Y VGND VGND VPWR VPWR _11903_/A sky130_fd_sc_hd__o21ai_1
X_12882_ _12853_/A _12853_/B _12853_/Y VGND VGND VPWR VPWR _12882_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14621_ _15341_/A _14655_/B VGND VGND VPWR VPWR _14621_/Y sky130_fd_sc_hd__nor2_1
X_11833_ _15143_/A _11838_/B VGND VGND VPWR VPWR _11833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14552_/A _14515_/X VGND VGND VPWR VPWR _14552_/X sky130_fd_sc_hd__or2b_1
X_11764_ _11764_/A VGND VGND VPWR VPWR _11808_/B sky130_fd_sc_hd__inv_2
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _15196_/A _14519_/B VGND VGND VPWR VPWR _14544_/A sky130_fd_sc_hd__and2_1
X_10715_ _10647_/A _10714_/Y _10647_/A _10714_/Y VGND VGND VPWR VPWR _10716_/B sky130_fd_sc_hd__a2bb2o_1
X_13503_ _13503_/A _13503_/B VGND VGND VPWR VPWR _13503_/Y sky130_fd_sc_hd__nand2_1
X_11695_ _11612_/Y _11692_/Y _11694_/X VGND VGND VPWR VPWR _11695_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16222_ _16089_/A _16089_/B _16089_/Y VGND VGND VPWR VPWR _16224_/A sky130_fd_sc_hd__o21ai_1
X_13434_ _13360_/X _13433_/X _13360_/X _13433_/X VGND VGND VPWR VPWR _13434_/Y sky130_fd_sc_hd__a2bb2oi_1
X_10646_ _10590_/Y _10644_/Y _10645_/Y VGND VGND VPWR VPWR _10647_/A sky130_fd_sc_hd__o21ai_1
X_16153_ _16270_/B VGND VGND VPWR VPWR _16336_/A sky130_fd_sc_hd__buf_6
Xrebuffer5 rebuffer6/X VGND VGND VPWR VPWR rebuffer5/X sky130_fd_sc_hd__dlygate4sd1_1
X_13365_ _13387_/A _13363_/X _13364_/X VGND VGND VPWR VPWR _13365_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10577_ _13515_/A _10667_/B _13515_/A _10667_/B VGND VGND VPWR VPWR _10577_/X sky130_fd_sc_hd__a2bb2o_1
X_15104_ _15104_/A _15104_/B VGND VGND VPWR VPWR _15105_/B sky130_fd_sc_hd__or2_1
X_16084_ _16084_/A _16084_/B VGND VGND VPWR VPWR _16084_/Y sky130_fd_sc_hd__nand2_1
X_12316_ _12324_/A VGND VGND VPWR VPWR _15512_/A sky130_fd_sc_hd__clkbuf_2
X_13296_ _13296_/A VGND VGND VPWR VPWR _13296_/Y sky130_fd_sc_hd__inv_2
X_12247_ _14057_/A _12211_/B _12211_/Y _12246_/X VGND VGND VPWR VPWR _12247_/X sky130_fd_sc_hd__a2bb2o_1
X_15035_ _15073_/A _15033_/X _15034_/X VGND VGND VPWR VPWR _15035_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12178_ _12178_/A VGND VGND VPWR VPWR _12270_/B sky130_fd_sc_hd__inv_2
XFILLER_110_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11129_ _11128_/A _11128_/B _11128_/X _10954_/X VGND VGND VPWR VPWR _11129_/X sky130_fd_sc_hd__o22a_1
XFILLER_1_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15937_ _15890_/A _15890_/B _15890_/Y VGND VGND VPWR VPWR _15937_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15868_ _15896_/A _15896_/B VGND VGND VPWR VPWR _15868_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14819_ _14806_/A _14806_/B _14806_/X _14818_/X VGND VGND VPWR VPWR _14819_/X sky130_fd_sc_hd__o22a_1
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15799_ _15670_/X _15798_/Y _15670_/X _15798_/Y VGND VGND VPWR VPWR _16217_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08340_ _08338_/Y _08339_/A _08338_/A _08339_/Y _08304_/A VGND VGND VPWR VPWR _09213_/B
+ sky130_fd_sc_hd__o221a_1
X_08271_ input27/X VGND VGND VPWR VPWR _08272_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_20_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09725_ _09770_/A _09770_/B VGND VGND VPWR VPWR _09725_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09656_ _09984_/A _09656_/B VGND VGND VPWR VPWR _09656_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _09456_/B VGND VGND VPWR VPWR _08716_/B sky130_fd_sc_hd__inv_2
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09587_ _09513_/X _09586_/X _09513_/X _09586_/X VGND VGND VPWR VPWR _09989_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08538_ _08538_/A VGND VGND VPWR VPWR _08538_/Y sky130_fd_sc_hd__clkinvlp_2
X_08469_ input22/X input6/X VGND VGND VPWR VPWR _08469_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10500_ _10499_/A _10498_/Y _10499_/Y _10498_/A _09941_/A VGND VGND VPWR VPWR _12928_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11480_ _15107_/A VGND VGND VPWR VPWR _13544_/A sky130_fd_sc_hd__buf_1
XFILLER_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10431_ _12826_/A _10431_/B VGND VGND VPWR VPWR _10431_/X sky130_fd_sc_hd__or2_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13150_ _13202_/A _13202_/B VGND VGND VPWR VPWR _13150_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10362_ _10362_/A VGND VGND VPWR VPWR _10362_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13081_ _13018_/X _13080_/X _13018_/X _13080_/X VGND VGND VPWR VPWR _13109_/B sky130_fd_sc_hd__a2bb2o_1
X_12101_ _13702_/A _12162_/B _12100_/Y VGND VGND VPWR VPWR _12101_/Y sky130_fd_sc_hd__o21ai_1
X_10293_ _10212_/X _12705_/A _10212_/X _12705_/A VGND VGND VPWR VPWR _10335_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12032_ _13190_/A _12057_/B VGND VGND VPWR VPWR _12032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13983_ _13984_/A _13984_/B VGND VGND VPWR VPWR _13983_/X sky130_fd_sc_hd__and2_1
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15722_ _16119_/A VGND VGND VPWR VPWR _15817_/A sky130_fd_sc_hd__inv_2
X_12934_ _12934_/A _12934_/B VGND VGND VPWR VPWR _12934_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15653_ _16030_/A VGND VGND VPWR VPWR _15667_/B sky130_fd_sc_hd__inv_2
X_12865_ _15171_/A _12864_/B _12864_/Y VGND VGND VPWR VPWR _12865_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15584_ _14394_/X _15583_/Y _14394_/X _15583_/Y VGND VGND VPWR VPWR _15685_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14604_/A _14603_/X VGND VGND VPWR VPWR _14604_/X sky130_fd_sc_hd__or2b_1
X_12796_ _12859_/A _12859_/B VGND VGND VPWR VPWR _12796_/Y sky130_fd_sc_hd__nor2_1
X_11816_ _12772_/A _11851_/A VGND VGND VPWR VPWR _11816_/Y sky130_fd_sc_hd__nor2_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _15190_/A _14535_/B VGND VGND VPWR VPWR _14535_/X sky130_fd_sc_hd__or2_1
X_11747_ _11745_/A _11745_/B _11745_/X _11746_/Y VGND VGND VPWR VPWR _11760_/B sky130_fd_sc_hd__a22o_1
XFILLER_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16205_ _16205_/A _16205_/B VGND VGND VPWR VPWR _16255_/A sky130_fd_sc_hd__or2_1
X_14466_ _14466_/A _14466_/B VGND VGND VPWR VPWR _14466_/Y sky130_fd_sc_hd__nand2_1
X_11678_ _12680_/A VGND VGND VPWR VPWR _12428_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14397_ _15970_/A _14400_/B VGND VGND VPWR VPWR _14397_/X sky130_fd_sc_hd__and2_1
X_13417_ _14095_/A _13420_/B VGND VGND VPWR VPWR _13417_/Y sky130_fd_sc_hd__nor2_1
X_10629_ _11892_/A _10629_/B VGND VGND VPWR VPWR _10629_/Y sky130_fd_sc_hd__nor2_1
X_16136_ _16136_/A _16136_/B VGND VGND VPWR VPWR _16136_/X sky130_fd_sc_hd__or2_1
XFILLER_127_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13348_ _13348_/A _13348_/B VGND VGND VPWR VPWR _13348_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16067_ _16114_/A _16114_/B VGND VGND VPWR VPWR _16067_/X sky130_fd_sc_hd__and2_1
XFILLER_6_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13279_ _14726_/A _13279_/B VGND VGND VPWR VPWR _13279_/Y sky130_fd_sc_hd__nand2_1
X_15018_ _15036_/A _15036_/B VGND VGND VPWR VPWR _15070_/A sky130_fd_sc_hd__and2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09510_ _09496_/A _09496_/B _09496_/Y _09509_/X VGND VGND VPWR VPWR _09510_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09441_ _09429_/A _09429_/B _09429_/X _09440_/X VGND VGND VPWR VPWR _09441_/X sky130_fd_sc_hd__a22o_2
XFILLER_24_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09372_ _09355_/X _09371_/X _09355_/X _09371_/X VGND VGND VPWR VPWR _09373_/A sky130_fd_sc_hd__a2bb2o_1
X_08323_ _08323_/A VGND VGND VPWR VPWR _08323_/Y sky130_fd_sc_hd__inv_2
X_08254_ input17/X _08254_/B VGND VGND VPWR VPWR _08327_/A sky130_fd_sc_hd__nor2_1
XFILLER_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09708_ _09681_/A _09101_/A _08928_/A _09707_/Y VGND VGND VPWR VPWR _09709_/B sky130_fd_sc_hd__o22a_1
XFILLER_55_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10980_ _10980_/A VGND VGND VPWR VPWR _10980_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09639_ _09543_/X _09638_/Y _09543_/X _09638_/Y VGND VGND VPWR VPWR _10743_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12650_ _12651_/A _12651_/B VGND VGND VPWR VPWR _12650_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11601_ _11577_/Y _10122_/Y _10237_/X VGND VGND VPWR VPWR _11602_/B sky130_fd_sc_hd__o21a_1
X_14320_ _14334_/A _14320_/B VGND VGND VPWR VPWR _15960_/A sky130_fd_sc_hd__or2_1
X_12581_ _12581_/A VGND VGND VPWR VPWR _12581_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11532_ _11615_/A _11615_/B _11531_/X VGND VGND VPWR VPWR _11533_/A sky130_fd_sc_hd__o21ai_1
X_14251_ _14233_/Y _14249_/Y _14250_/Y VGND VGND VPWR VPWR _14252_/A sky130_fd_sc_hd__o21ai_1
XFILLER_11_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11463_ _08983_/X _11462_/X _08983_/X _11462_/X VGND VGND VPWR VPWR _11464_/B sky130_fd_sc_hd__a2bb2oi_2
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14182_ _14281_/A _14182_/B VGND VGND VPWR VPWR _15857_/A sky130_fd_sc_hd__or2_1
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13202_ _13202_/A _13202_/B VGND VGND VPWR VPWR _13202_/Y sky130_fd_sc_hd__nand2_1
X_10414_ _10357_/X _10413_/X _10357_/X _10413_/X VGND VGND VPWR VPWR _10431_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11394_ _14102_/A VGND VGND VPWR VPWR _12346_/A sky130_fd_sc_hd__inv_2
X_13133_ _13133_/A VGND VGND VPWR VPWR _13966_/A sky130_fd_sc_hd__inv_2
XFILLER_124_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10345_ _10421_/A VGND VGND VPWR VPWR _10424_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_3_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13064_ _13768_/A VGND VGND VPWR VPWR _15249_/A sky130_fd_sc_hd__buf_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10276_ _10228_/A _10228_/B _10228_/Y VGND VGND VPWR VPWR _10277_/A sky130_fd_sc_hd__a21oi_2
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ _11979_/X _12014_/Y _11979_/X _12014_/Y VGND VGND VPWR VPWR _12065_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13966_ _13966_/A _13967_/B VGND VGND VPWR VPWR _13968_/A sky130_fd_sc_hd__and2_1
X_15705_ _15697_/X _15704_/Y _15697_/X _15704_/Y VGND VGND VPWR VPWR _15823_/B sky130_fd_sc_hd__a2bb2o_1
X_13897_ _13897_/A VGND VGND VPWR VPWR _15414_/A sky130_fd_sc_hd__buf_1
X_12917_ _12917_/A VGND VGND VPWR VPWR _12917_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15636_ _14347_/X _15636_/B VGND VGND VPWR VPWR _15636_/Y sky130_fd_sc_hd__nand2b_1
X_12848_ _12814_/Y _12846_/X _12847_/Y VGND VGND VPWR VPWR _12848_/X sky130_fd_sc_hd__o21a_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ _15565_/X _15566_/X _15565_/X _15566_/X VGND VGND VPWR VPWR _15567_/Y sky130_fd_sc_hd__a2bb2oi_1
X_12779_ _12739_/Y _12777_/X _12778_/Y VGND VGND VPWR VPWR _12779_/X sky130_fd_sc_hd__o21a_1
X_15498_ _15446_/A _15446_/B _15446_/A _15446_/B VGND VGND VPWR VPWR _15498_/X sky130_fd_sc_hd__a2bb2o_1
X_14518_ _14548_/A _14516_/X _14517_/X VGND VGND VPWR VPWR _14518_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14449_ _14432_/X _14448_/X _14432_/X _14448_/X VGND VGND VPWR VPWR _14462_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16119_ _16119_/A _16119_/B VGND VGND VPWR VPWR _16119_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09990_ _09990_/A _09990_/B VGND VGND VPWR VPWR _09990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08941_ _08678_/A _08940_/X _08678_/A _08940_/X VGND VGND VPWR VPWR _11407_/A sky130_fd_sc_hd__a2bb2o_1
X_08872_ _08693_/X _08871_/Y _08693_/X _08871_/Y VGND VGND VPWR VPWR _08984_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09424_ _09424_/A _09424_/B VGND VGND VPWR VPWR _09424_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09355_ _08690_/A _09860_/A _09352_/Y _09354_/X VGND VGND VPWR VPWR _09355_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08306_ input22/X _08306_/B VGND VGND VPWR VPWR _08307_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09286_ _09254_/Y _08954_/Y _09254_/Y _08954_/Y VGND VGND VPWR VPWR _10245_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08237_ _08237_/A input23/X VGND VGND VPWR VPWR _08238_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10130_ _10130_/A _10130_/B VGND VGND VPWR VPWR _10131_/B sky130_fd_sc_hd__or2_1
XFILLER_88_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10061_ _10061_/A _10061_/B VGND VGND VPWR VPWR _10061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13820_ _14626_/A _13845_/B VGND VGND VPWR VPWR _13820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13751_ _11961_/X _13750_/X _11961_/X _13750_/X VGND VGND VPWR VPWR _13752_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10963_ _12082_/A VGND VGND VPWR VPWR _11999_/A sky130_fd_sc_hd__inv_2
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16470_ _08229_/A _16470_/D VGND VGND VPWR VPWR _16470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12702_ _12702_/A VGND VGND VPWR VPWR _12704_/A sky130_fd_sc_hd__buf_1
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15421_ _15359_/X _15419_/X _15435_/B VGND VGND VPWR VPWR _15421_/Y sky130_fd_sc_hd__o21ai_1
X_10894_ _12039_/A _10894_/B VGND VGND VPWR VPWR _10894_/Y sky130_fd_sc_hd__nor2_1
X_13682_ _12921_/A _13681_/X _12921_/A _13681_/X VGND VGND VPWR VPWR _13683_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12633_ _14189_/A _12631_/X _12632_/X VGND VGND VPWR VPWR _12633_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12564_ _12561_/Y _12563_/Y _12561_/A _12563_/A _12503_/A VGND VGND VPWR VPWR _12626_/B
+ sky130_fd_sc_hd__o221a_1
X_15352_ _15296_/X _15350_/X _15360_/B VGND VGND VPWR VPWR _15352_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14303_ _15906_/A _14277_/B _14277_/Y VGND VGND VPWR VPWR _14303_/Y sky130_fd_sc_hd__o21ai_1
X_15283_ _14833_/A _15237_/B _15237_/Y _15282_/X VGND VGND VPWR VPWR _15283_/X sky130_fd_sc_hd__a2bb2o_1
X_11515_ _11629_/A VGND VGND VPWR VPWR _13495_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14234_ _14234_/A _14234_/B VGND VGND VPWR VPWR _15839_/A sky130_fd_sc_hd__nor2_1
X_12495_ _12410_/A _12410_/B _12410_/Y _12412_/A VGND VGND VPWR VPWR _12495_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_125_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11446_ _14027_/A _11219_/B _11219_/Y VGND VGND VPWR VPWR _11446_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14165_ _15974_/A _14165_/B VGND VGND VPWR VPWR _14166_/B sky130_fd_sc_hd__or2_1
X_11377_ _14057_/A _11197_/B _11197_/Y VGND VGND VPWR VPWR _11377_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14096_ _14092_/Y _14094_/Y _14095_/Y VGND VGND VPWR VPWR _14100_/B sky130_fd_sc_hd__o21ai_1
X_13116_ _13067_/Y _13114_/X _13115_/Y VGND VGND VPWR VPWR _13116_/X sky130_fd_sc_hd__o21a_1
X_10328_ _13527_/A _10328_/B VGND VGND VPWR VPWR _10328_/X sky130_fd_sc_hd__and2_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _15237_/A _13123_/B VGND VGND VPWR VPWR _13047_/Y sky130_fd_sc_hd__nor2_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10259_ _09262_/B _10242_/B _10242_/X _10829_/A VGND VGND VPWR VPWR _10983_/A sky130_fd_sc_hd__a22o_1
XFILLER_120_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14998_ _11734_/A _11733_/Y _11727_/Y _14997_/X VGND VGND VPWR VPWR _14998_/X sky130_fd_sc_hd__o22a_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13949_ _15408_/A _13949_/B VGND VGND VPWR VPWR _13949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15619_ _16038_/A VGND VGND VPWR VPWR _15675_/A sky130_fd_sc_hd__inv_2
XFILLER_62_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09140_ _09140_/A VGND VGND VPWR VPWR _09140_/Y sky130_fd_sc_hd__inv_2
X_09071_ _10018_/B _09071_/B VGND VGND VPWR VPWR _09072_/B sky130_fd_sc_hd__or2_1
XFILLER_30_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09973_ _09963_/Y _09972_/Y _09960_/Y VGND VGND VPWR VPWR _09975_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08924_ _09541_/A _10098_/B _08678_/A VGND VGND VPWR VPWR _08932_/B sky130_fd_sc_hd__o21ai_1
XFILLER_130_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08855_ _09503_/A _09041_/B VGND VGND VPWR VPWR _08855_/Y sky130_fd_sc_hd__nor2_1
X_08786_ _09470_/A _08786_/B VGND VGND VPWR VPWR _08786_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09407_ _09407_/A _09407_/B VGND VGND VPWR VPWR _09407_/X sky130_fd_sc_hd__or2_1
X_09338_ _09448_/A _09338_/B VGND VGND VPWR VPWR _09338_/X sky130_fd_sc_hd__or2_1
XFILLER_40_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11300_ _11300_/A _11300_/B VGND VGND VPWR VPWR _11300_/Y sky130_fd_sc_hd__nor2_1
X_09269_ _08597_/A _09856_/A _09216_/A VGND VGND VPWR VPWR _09269_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12280_ _12371_/B _12279_/Y _12371_/B _12279_/Y VGND VGND VPWR VPWR _12369_/B sky130_fd_sc_hd__o2bb2a_1
X_11231_ _14035_/A _11231_/B VGND VGND VPWR VPWR _11231_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11162_ _12261_/A _11304_/B _12261_/A _11304_/B VGND VGND VPWR VPWR _11162_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10113_ _10113_/A _10113_/B VGND VGND VPWR VPWR _10114_/A sky130_fd_sc_hd__or2_1
XFILLER_121_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15970_ _15970_/A _15970_/B VGND VGND VPWR VPWR _15970_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11093_ _11195_/A _11091_/X _11092_/X VGND VGND VPWR VPWR _11093_/X sky130_fd_sc_hd__o21a_1
X_14921_ _14879_/Y _14919_/X _14920_/Y VGND VGND VPWR VPWR _14921_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10044_ _10044_/A _10044_/B VGND VGND VPWR VPWR _10044_/Y sky130_fd_sc_hd__nor2_1
X_14852_ _14953_/A _14953_/B _14851_/Y VGND VGND VPWR VPWR _14852_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13803_ _13803_/A _13772_/X VGND VGND VPWR VPWR _13803_/X sky130_fd_sc_hd__or2b_1
XFILLER_29_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14783_ _15449_/A VGND VGND VPWR VPWR _14786_/A sky130_fd_sc_hd__buf_1
XFILLER_91_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11995_ _10682_/A _11925_/A _10814_/B _11994_/Y VGND VGND VPWR VPWR _11996_/A sky130_fd_sc_hd__o22a_1
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13734_ _13766_/A _13766_/B VGND VGND VPWR VPWR _13812_/A sky130_fd_sc_hd__and2_1
X_10946_ _13640_/A _10946_/B VGND VGND VPWR VPWR _10946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16453_ _16349_/X _16406_/A _16409_/A VGND VGND VPWR VPWR _16454_/B sky130_fd_sc_hd__o21a_1
X_10877_ _10775_/X _10876_/Y _10775_/X _10876_/Y VGND VGND VPWR VPWR _10878_/B sky130_fd_sc_hd__o2bb2a_1
X_13665_ _13627_/A _13664_/Y _13627_/A _13664_/Y VGND VGND VPWR VPWR _13694_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16384_ _16160_/A _16384_/B VGND VGND VPWR VPWR _16395_/A sky130_fd_sc_hd__nand2b_1
X_12616_ _14234_/A _14234_/B VGND VGND VPWR VPWR _12617_/A sky130_fd_sc_hd__nand2_1
X_15404_ _15404_/A _15404_/B VGND VGND VPWR VPWR _15404_/X sky130_fd_sc_hd__or2_1
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15335_ _15335_/A _15335_/B VGND VGND VPWR VPWR _15335_/X sky130_fd_sc_hd__or2_1
X_13596_ _13559_/A _13559_/B _13560_/A VGND VGND VPWR VPWR _13596_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12547_ _15540_/A VGND VGND VPWR VPWR _14916_/A sky130_fd_sc_hd__buf_1
X_12478_ _13462_/A _12480_/B VGND VGND VPWR VPWR _12478_/Y sky130_fd_sc_hd__nor2_1
X_15266_ _15217_/X _15265_/Y _15217_/X _15265_/Y VGND VGND VPWR VPWR _15272_/B sky130_fd_sc_hd__a2bb2o_1
XANTENNA_3 _08656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14217_ _14094_/Y _14216_/X _14094_/Y _14216_/X VGND VGND VPWR VPWR _14218_/B sky130_fd_sc_hd__a2bb2oi_1
X_11429_ _14038_/A _11238_/B _11238_/Y VGND VGND VPWR VPWR _11429_/Y sky130_fd_sc_hd__o21ai_1
X_15197_ _15131_/A _15131_/B _15131_/Y VGND VGND VPWR VPWR _15197_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14148_ _14148_/A _14148_/B VGND VGND VPWR VPWR _14148_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ _14815_/A _14047_/B _14047_/Y VGND VGND VPWR VPWR _14079_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08640_ _09459_/B VGND VGND VPWR VPWR _08719_/B sky130_fd_sc_hd__inv_2
XFILLER_94_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer26 _08395_/A VGND VGND VPWR VPWR _08666_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer15 rebuffer16/X VGND VGND VPWR VPWR rebuffer15/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer59 _11723_/B VGND VGND VPWR VPWR _11716_/B sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer48 _08375_/X VGND VGND VPWR VPWR _08454_/A sky130_fd_sc_hd__dlygate4sd1_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08571_ _08571_/A VGND VGND VPWR VPWR _10116_/B sky130_fd_sc_hd__inv_2
Xrebuffer37 _09748_/A VGND VGND VPWR VPWR _09750_/B sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_22_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09123_ _09703_/A _09123_/B VGND VGND VPWR VPWR _09123_/Y sky130_fd_sc_hd__nand2_1
X_09054_ _09054_/A VGND VGND VPWR VPWR _09054_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09956_ _09955_/A _09955_/B _09954_/Y _09955_/X VGND VGND VPWR VPWR _09958_/B sky130_fd_sc_hd__o22ai_2
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09887_/A _09887_/B VGND VGND VPWR VPWR _09888_/B sky130_fd_sc_hd__or2_1
X_08907_ _08972_/A _08972_/B VGND VGND VPWR VPWR _08907_/X sky130_fd_sc_hd__and2_1
XFILLER_85_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _08718_/A _09462_/B _08718_/Y VGND VGND VPWR VPWR _08839_/A sky130_fd_sc_hd__a21oi_2
XFILLER_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08769_ _10010_/A VGND VGND VPWR VPWR _08770_/A sky130_fd_sc_hd__buf_1
XFILLER_122_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11780_ _12766_/A _11780_/B VGND VGND VPWR VPWR _11780_/Y sky130_fd_sc_hd__nor2_1
X_10800_ _09262_/A _09262_/B _09262_/X VGND VGND VPWR VPWR _10801_/B sky130_fd_sc_hd__a21boi_1
X_10731_ _13692_/A _10642_/B _10642_/Y VGND VGND VPWR VPWR _10731_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13450_ _13374_/Y _13448_/X _13449_/Y VGND VGND VPWR VPWR _13450_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12401_ _12399_/X _12401_/B VGND VGND VPWR VPWR _12401_/Y sky130_fd_sc_hd__nand2b_1
X_10662_ _10545_/X _10661_/B _10661_/X _10541_/X VGND VGND VPWR VPWR _10662_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13381_ _13381_/A _13368_/X VGND VGND VPWR VPWR _13381_/X sky130_fd_sc_hd__or2b_1
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10593_ _09971_/Y _10592_/A _09971_/A _10592_/Y _09797_/A VGND VGND VPWR VPWR _11904_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_126_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12332_ _12591_/A _12590_/A _12331_/X VGND VGND VPWR VPWR _12336_/B sky130_fd_sc_hd__o21ai_2
X_15120_ _15063_/A _15063_/B _15063_/Y VGND VGND VPWR VPWR _15120_/Y sky130_fd_sc_hd__o21ai_1
X_12263_ _12263_/A _12263_/B VGND VGND VPWR VPWR _12263_/X sky130_fd_sc_hd__or2_1
X_15051_ _15051_/A _15051_/B VGND VGND VPWR VPWR _15052_/B sky130_fd_sc_hd__or2_1
XFILLER_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14002_ _14067_/A _14067_/B VGND VGND VPWR VPWR _14002_/X sky130_fd_sc_hd__and2_1
X_11214_ _11214_/A _11220_/B VGND VGND VPWR VPWR _13334_/A sky130_fd_sc_hd__or2_1
XFILLER_134_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12194_ _12257_/A _12193_/Y _12257_/A _12193_/Y VGND VGND VPWR VPWR _12254_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11145_ _11145_/A VGND VGND VPWR VPWR _12270_/A sky130_fd_sc_hd__inv_2
X_15953_ _15939_/X _15951_/X _16017_/B VGND VGND VPWR VPWR _15953_/X sky130_fd_sc_hd__o21a_1
X_11076_ _13935_/A _12234_/B _11074_/X _11248_/A VGND VGND VPWR VPWR _11076_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14904_ _14904_/A _14904_/B VGND VGND VPWR VPWR _14904_/Y sky130_fd_sc_hd__nor2_1
X_10027_ _09452_/A _08786_/B _10044_/B _10026_/X VGND VGND VPWR VPWR _10027_/X sky130_fd_sc_hd__o22a_1
X_15884_ _14242_/A _15839_/B _14236_/A _14370_/X _14242_/B VGND VGND VPWR VPWR _15885_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_91_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14835_ _14748_/X _14762_/A _14761_/X VGND VGND VPWR VPWR _14835_/X sky130_fd_sc_hd__o21a_1
X_14766_ _14746_/X _14765_/Y _14746_/X _14765_/Y VGND VGND VPWR VPWR _14830_/B sky130_fd_sc_hd__a2bb2o_1
X_11978_ _13063_/A _11978_/B VGND VGND VPWR VPWR _11978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13717_ _13777_/A _13716_/Y _13777_/A _13716_/Y VGND VGND VPWR VPWR _13719_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10929_ _10929_/A VGND VGND VPWR VPWR _11586_/A sky130_fd_sc_hd__clkbuf_2
X_14697_ _14656_/X _14696_/Y _14656_/X _14696_/Y VGND VGND VPWR VPWR _14734_/B sky130_fd_sc_hd__a2bb2o_1
X_16436_ _16460_/Q _16459_/Q _16465_/Q _16435_/X _16437_/D VGND VGND VPWR VPWR _16436_/X
+ sky130_fd_sc_hd__o41a_1
X_13648_ _13648_/A _13648_/B VGND VGND VPWR VPWR _13708_/A sky130_fd_sc_hd__nand2_1
X_16367_ _16325_/X _16366_/Y _16325_/X _16366_/Y VGND VGND VPWR VPWR _16407_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13579_ _12849_/A _13551_/B _13552_/Y _13578_/X VGND VGND VPWR VPWR _13579_/X sky130_fd_sc_hd__o22a_1
X_16298_ _16259_/X _16297_/Y _16259_/X _16297_/Y VGND VGND VPWR VPWR _16326_/B sky130_fd_sc_hd__o2bb2a_1
X_15318_ _14577_/A _15261_/B _15261_/Y VGND VGND VPWR VPWR _15318_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15249_ _15249_/A _15249_/B VGND VGND VPWR VPWR _15249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09810_ _09458_/Y _09809_/X _09462_/X VGND VGND VPWR VPWR _09810_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09741_ _08535_/A _09743_/B _08535_/A _09743_/B VGND VGND VPWR VPWR _09742_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09672_ _09672_/A VGND VGND VPWR VPWR _10933_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08623_ _08623_/A _10112_/B VGND VGND VPWR VPWR _08624_/A sky130_fd_sc_hd__or2_1
XFILLER_27_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _08554_/A VGND VGND VPWR VPWR _10011_/A sky130_fd_sc_hd__buf_1
XFILLER_63_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08485_ _08272_/A _08363_/B _08479_/Y _08625_/A VGND VGND VPWR VPWR _08612_/A sky130_fd_sc_hd__o22a_1
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09106_ _09407_/A _09104_/B _09104_/X _09105_/X VGND VGND VPWR VPWR _09107_/B sky130_fd_sc_hd__o22a_1
X_09037_ _09531_/B _09037_/B VGND VGND VPWR VPWR _09038_/B sky130_fd_sc_hd__or2_1
XFILLER_123_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09939_ _09935_/Y _09938_/X _09935_/Y _09938_/X VGND VGND VPWR VPWR _11595_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12950_ _12868_/Y _12947_/X _12949_/Y VGND VGND VPWR VPWR _12950_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11901_ _12992_/A _11901_/B VGND VGND VPWR VPWR _11901_/Y sky130_fd_sc_hd__nand2_1
X_12881_ _12940_/A VGND VGND VPWR VPWR _14531_/A sky130_fd_sc_hd__buf_1
XFILLER_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14620_ _14582_/X _14619_/Y _14582_/X _14619_/Y VGND VGND VPWR VPWR _14655_/B sky130_fd_sc_hd__a2bb2o_1
X_11832_ _11796_/X _11831_/X _11796_/X _11831_/X VGND VGND VPWR VPWR _11838_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _15258_/A VGND VGND VPWR VPWR _14579_/A sky130_fd_sc_hd__buf_1
XFILLER_73_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _10303_/A _11750_/A _10369_/B _11762_/Y VGND VGND VPWR VPWR _11764_/A sky130_fd_sc_hd__o22a_1
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14467_/X _14481_/Y _14467_/X _14481_/Y VGND VGND VPWR VPWR _14519_/B sky130_fd_sc_hd__a2bb2o_1
X_10714_ _13696_/A _10648_/B _10648_/Y VGND VGND VPWR VPWR _10714_/Y sky130_fd_sc_hd__o21ai_1
X_13502_ _11158_/X _13489_/X _11158_/X _13489_/X VGND VGND VPWR VPWR _13503_/B sky130_fd_sc_hd__o2bb2a_1
X_11694_ _12426_/A _11694_/B VGND VGND VPWR VPWR _11694_/X sky130_fd_sc_hd__or2_1
X_16221_ _16253_/A _16320_/A VGND VGND VPWR VPWR _16221_/Y sky130_fd_sc_hd__nor2_1
X_13433_ _13331_/A _13331_/B _13331_/A _13331_/B VGND VGND VPWR VPWR _13433_/X sky130_fd_sc_hd__a2bb2o_1
X_10645_ _11907_/A _10645_/B VGND VGND VPWR VPWR _10645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16152_ _16160_/A _16152_/B VGND VGND VPWR VPWR _16270_/B sky130_fd_sc_hd__or2_1
X_13364_ _13364_/A _13364_/B VGND VGND VPWR VPWR _13364_/X sky130_fd_sc_hd__or2_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12315_ _14083_/A VGND VGND VPWR VPWR _12324_/A sky130_fd_sc_hd__inv_2
X_15103_ _15104_/A _15104_/B VGND VGND VPWR VPWR _15103_/X sky130_fd_sc_hd__and2_1
X_10576_ _10555_/X _10575_/X _10555_/X _10575_/X VGND VGND VPWR VPWR _10667_/B sky130_fd_sc_hd__a2bb2o_1
Xrebuffer6 rebuffer7/X VGND VGND VPWR VPWR rebuffer6/X sky130_fd_sc_hd__dlygate4sd1_1
X_16083_ _15781_/A _15766_/A _15784_/B VGND VGND VPWR VPWR _16233_/A sky130_fd_sc_hd__o21ai_2
XFILLER_108_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13295_ _13235_/Y _13293_/Y _13294_/Y VGND VGND VPWR VPWR _13296_/A sky130_fd_sc_hd__o21ai_1
XFILLER_108_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12246_ _14055_/A _12214_/B _12214_/Y _12245_/X VGND VGND VPWR VPWR _12246_/X sky130_fd_sc_hd__a2bb2o_1
X_15034_ _15034_/A _15034_/B VGND VGND VPWR VPWR _15034_/X sky130_fd_sc_hd__or2_1
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12177_ _10972_/A _12086_/A _11140_/B _12176_/Y VGND VGND VPWR VPWR _12178_/A sky130_fd_sc_hd__o22a_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11128_ _11128_/A _11128_/B VGND VGND VPWR VPWR _11128_/X sky130_fd_sc_hd__and2_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15936_ _15954_/A _15954_/B VGND VGND VPWR VPWR _15936_/X sky130_fd_sc_hd__and2_1
X_11059_ _12139_/A _11078_/B VGND VGND VPWR VPWR _11242_/A sky130_fd_sc_hd__and2_1
XFILLER_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15867_ _14201_/X _15845_/X _14201_/X _15845_/X VGND VGND VPWR VPWR _15896_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14818_ _14809_/A _14809_/B _14809_/Y _14817_/X VGND VGND VPWR VPWR _14818_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15798_ _15671_/A _15671_/B _15671_/Y VGND VGND VPWR VPWR _15798_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14749_ _14749_/A VGND VGND VPWR VPWR _15181_/A sky130_fd_sc_hd__buf_1
X_08270_ input11/X VGND VGND VPWR VPWR _08363_/B sky130_fd_sc_hd__clkinvlp_2
X_16419_ _16474_/Q _16419_/B VGND VGND VPWR VPWR _16429_/B sky130_fd_sc_hd__or2_1
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09724_ _09970_/A _09722_/Y _09723_/Y VGND VGND VPWR VPWR _09770_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09655_ _09609_/Y _09653_/X _09654_/Y VGND VGND VPWR VPWR _09655_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08606_ _08605_/X _08417_/Y _08605_/X _08417_/Y VGND VGND VPWR VPWR _08609_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09586_ _09488_/A _09488_/B _09488_/Y VGND VGND VPWR VPWR _09586_/X sky130_fd_sc_hd__a21o_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08692_/A _10119_/B VGND VGND VPWR VPWR _08876_/A sky130_fd_sc_hd__nor2_1
X_08468_ _08505_/B _08464_/Y _08704_/B VGND VGND VPWR VPWR _08468_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_23_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10430_ _12827_/A _10429_/B _10428_/X _10429_/X VGND VGND VPWR VPWR _10430_/X sky130_fd_sc_hd__o22a_1
X_08399_ _08399_/A _08399_/B VGND VGND VPWR VPWR _08662_/B sky130_fd_sc_hd__or2_1
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10361_ _09975_/A _09975_/B _09975_/Y VGND VGND VPWR VPWR _10362_/A sky130_fd_sc_hd__o21ai_1
XFILLER_124_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13080_ _13080_/A _13019_/X VGND VGND VPWR VPWR _13080_/X sky130_fd_sc_hd__or2b_1
X_12100_ _12162_/A _12162_/B VGND VGND VPWR VPWR _12100_/Y sky130_fd_sc_hd__nand2_1
X_10292_ _10213_/A _10213_/B _10213_/Y VGND VGND VPWR VPWR _12705_/A sky130_fd_sc_hd__o21ai_2
X_12031_ _11971_/X _12030_/Y _11971_/X _12030_/Y VGND VGND VPWR VPWR _12057_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13982_ _13979_/Y _13981_/X _13979_/Y _13981_/X VGND VGND VPWR VPWR _13984_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15721_ _15728_/A _15721_/B VGND VGND VPWR VPWR _16119_/A sky130_fd_sc_hd__or2_1
X_12933_ _12900_/Y _12931_/X _12932_/Y VGND VGND VPWR VPWR _12933_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15652_ _15651_/A _15650_/Y _15651_/Y _15650_/A _15571_/A VGND VGND VPWR VPWR _16030_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_73_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12864_ _12864_/A _12864_/B VGND VGND VPWR VPWR _12864_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15583_ _14305_/X _15583_/B VGND VGND VPWR VPWR _15583_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _15187_/A _14603_/B VGND VGND VPWR VPWR _14603_/X sky130_fd_sc_hd__or2_1
XFILLER_61_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12795_ _12783_/X _12794_/Y _12783_/X _12794_/Y VGND VGND VPWR VPWR _12859_/B sky130_fd_sc_hd__a2bb2o_1
X_11815_ _11855_/B _11814_/Y _11855_/B _11814_/Y VGND VGND VPWR VPWR _11851_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _15190_/A _14535_/B VGND VGND VPWR VPWR _14536_/A sky130_fd_sc_hd__and2_1
X_11746_ _11746_/A VGND VGND VPWR VPWR _11746_/Y sky130_fd_sc_hd__inv_4
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16204_ _16098_/X _16203_/X _16098_/X _16203_/X VGND VGND VPWR VPWR _16205_/B sky130_fd_sc_hd__o2bb2a_1
X_11677_ _11674_/X _12644_/A _12643_/B VGND VGND VPWR VPWR _11677_/Y sky130_fd_sc_hd__o21ai_1
X_14465_ _14447_/Y _14463_/X _14464_/Y VGND VGND VPWR VPWR _14465_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14396_ _14305_/X _14394_/X _15583_/B VGND VGND VPWR VPWR _14400_/B sky130_fd_sc_hd__o21ai_1
X_13416_ _13412_/X _13414_/Y _14350_/B VGND VGND VPWR VPWR _13420_/B sky130_fd_sc_hd__o21ai_2
X_10628_ _11889_/A _15212_/B VGND VGND VPWR VPWR _10766_/A sky130_fd_sc_hd__or2_1
XFILLER_127_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16135_ _16388_/A _16135_/B VGND VGND VPWR VPWR _16136_/B sky130_fd_sc_hd__or2_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13347_ _13273_/X _13346_/Y _13273_/X _13346_/Y VGND VGND VPWR VPWR _13348_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10559_ _09088_/A _10558_/X _09088_/A _10558_/X VGND VGND VPWR VPWR _11207_/A sky130_fd_sc_hd__a2bb2o_2
X_16066_ _16045_/X _16065_/Y _16045_/X _16065_/Y VGND VGND VPWR VPWR _16114_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13278_ _13278_/A VGND VGND VPWR VPWR _13278_/Y sky130_fd_sc_hd__inv_2
X_12229_ _12229_/A _12229_/B VGND VGND VPWR VPWR _12229_/Y sky130_fd_sc_hd__nand2_1
X_15017_ _11814_/Y _15001_/X _11814_/Y _15001_/X VGND VGND VPWR VPWR _15036_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15919_ _15902_/A _15902_/B _15902_/Y VGND VGND VPWR VPWR _15919_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09440_ _09430_/A _09430_/B _09430_/X _09439_/X VGND VGND VPWR VPWR _09440_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09371_ _09474_/B _09861_/A _09350_/A VGND VGND VPWR VPWR _09371_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08322_ _08322_/A _08322_/B VGND VGND VPWR VPWR _08323_/A sky130_fd_sc_hd__or2_1
XFILLER_33_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08253_ input33/X VGND VGND VPWR VPWR _08254_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_32_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09707_ _09707_/A _09707_/B VGND VGND VPWR VPWR _09707_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09638_ _09539_/A _09539_/B _09539_/X VGND VGND VPWR VPWR _09638_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09569_ _09569_/A _09569_/B VGND VGND VPWR VPWR _09569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12580_ _12576_/Y _12579_/Y _12576_/A _12579_/A _11709_/A VGND VGND VPWR VPWR _12622_/A
+ sky130_fd_sc_hd__o221a_1
X_11600_ _15163_/A VGND VGND VPWR VPWR _12413_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_24_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11531_ _11531_/A _11531_/B VGND VGND VPWR VPWR _11531_/X sky130_fd_sc_hd__or2_1
XFILLER_11_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14250_ _15881_/A _14250_/B VGND VGND VPWR VPWR _14250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11462_ _08875_/X _11462_/B VGND VGND VPWR VPWR _11462_/X sky130_fd_sc_hd__and2b_1
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14181_ _14121_/X _14180_/Y _14121_/X _14180_/Y VGND VGND VPWR VPWR _14182_/B sky130_fd_sc_hd__a2bb2oi_1
X_11393_ _11393_/A _11393_/B VGND VGND VPWR VPWR _14102_/A sky130_fd_sc_hd__or2_1
X_13201_ _13153_/Y _13199_/X _13200_/Y VGND VGND VPWR VPWR _13201_/X sky130_fd_sc_hd__o21a_1
X_10413_ _13529_/A _10338_/B _11787_/A _10338_/B VGND VGND VPWR VPWR _10413_/X sky130_fd_sc_hd__a2bb2o_1
X_13132_ _13132_/A VGND VGND VPWR VPWR _14067_/A sky130_fd_sc_hd__inv_2
X_10344_ _12606_/A _10344_/B VGND VGND VPWR VPWR _10421_/A sky130_fd_sc_hd__or2_1
XFILLER_3_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13063_ _13063_/A VGND VGND VPWR VPWR _13768_/A sky130_fd_sc_hd__inv_2
X_10275_ _11727_/A VGND VGND VPWR VPWR _12707_/A sky130_fd_sc_hd__buf_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ _12068_/A _12068_/B _12013_/Y VGND VGND VPWR VPWR _12014_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13965_ _13542_/X _13964_/X _13542_/X _13964_/X VGND VGND VPWR VPWR _13967_/B sky130_fd_sc_hd__a2bb2o_1
X_15704_ _15991_/A _15825_/B _15703_/Y VGND VGND VPWR VPWR _15704_/Y sky130_fd_sc_hd__o21ai_1
X_13896_ _15416_/A _13957_/B VGND VGND VPWR VPWR _13896_/Y sky130_fd_sc_hd__nor2_1
X_12916_ _12915_/A _12915_/B _12915_/Y VGND VGND VPWR VPWR _12916_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ _16034_/A VGND VGND VPWR VPWR _15671_/A sky130_fd_sc_hd__inv_2
X_12847_ _12847_/A _12847_/B VGND VGND VPWR VPWR _12847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _15289_/A _15289_/B _15289_/Y _15354_/X VGND VGND VPWR VPWR _15566_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12778_ _12778_/A _12778_/B VGND VGND VPWR VPWR _12778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15497_ _15548_/A _15548_/B VGND VGND VPWR VPWR _15497_/X sky130_fd_sc_hd__and2_1
X_14517_ _15199_/A _14517_/B VGND VGND VPWR VPWR _14517_/X sky130_fd_sc_hd__or2_1
X_11729_ _11734_/B _11728_/Y _11734_/B _11728_/Y VGND VGND VPWR VPWR _11787_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14448_ _14424_/A _14424_/B _14424_/Y VGND VGND VPWR VPWR _14448_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14379_ _14379_/A _15950_/A VGND VGND VPWR VPWR _15644_/B sky130_fd_sc_hd__or2_1
X_16118_ _16050_/X _16117_/Y _16050_/X _16117_/Y VGND VGND VPWR VPWR _16147_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16049_ _15966_/A _15966_/B _15966_/Y VGND VGND VPWR VPWR _16049_/Y sky130_fd_sc_hd__o21ai_1
X_08940_ _08679_/A _08679_/B _08679_/A _08679_/B VGND VGND VPWR VPWR _08940_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08871_ _08871_/A _08871_/B VGND VGND VPWR VPWR _08871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09423_ _09769_/A _09424_/B VGND VGND VPWR VPWR _09423_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09354_ _08688_/A _09859_/A _09353_/Y _09318_/X VGND VGND VPWR VPWR _09354_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08305_ _08239_/Y _08296_/A _08239_/A _08296_/Y _08304_/X VGND VGND VPWR VPWR _08505_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09285_ _09285_/A VGND VGND VPWR VPWR _09285_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08236_ input7/X VGND VGND VPWR VPWR _08237_/A sky130_fd_sc_hd__inv_2
XFILLER_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10060_ _10059_/A _10059_/B _10216_/A _10059_/Y VGND VGND VPWR VPWR _10063_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13750_ _13683_/A _13683_/B _13683_/A _13683_/B VGND VGND VPWR VPWR _13750_/X sky130_fd_sc_hd__a2bb2o_1
X_10962_ _10964_/A VGND VGND VPWR VPWR _10962_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12701_ _12701_/A _12701_/B VGND VGND VPWR VPWR _12701_/Y sky130_fd_sc_hd__nor2_1
X_15420_ _15420_/A _15420_/B VGND VGND VPWR VPWR _15435_/B sky130_fd_sc_hd__or2_1
X_10893_ _10773_/X _10892_/Y _10773_/X _10892_/Y VGND VGND VPWR VPWR _10894_/B sky130_fd_sc_hd__a2bb2o_1
X_13681_ _13005_/A _13611_/A _13609_/Y _13611_/Y VGND VGND VPWR VPWR _13681_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12632_ _12632_/A _12632_/B VGND VGND VPWR VPWR _12632_/X sky130_fd_sc_hd__or2_1
XFILLER_31_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12563_ _12563_/A VGND VGND VPWR VPWR _12563_/Y sky130_fd_sc_hd__inv_2
X_15351_ _15351_/A _15351_/B VGND VGND VPWR VPWR _15360_/B sky130_fd_sc_hd__or2_1
X_14302_ _14308_/A _14302_/B VGND VGND VPWR VPWR _15966_/A sky130_fd_sc_hd__or2_1
X_12494_ _12496_/A _12496_/B VGND VGND VPWR VPWR _12494_/Y sky130_fd_sc_hd__nor2_1
X_15282_ _14745_/A _15240_/B _15240_/Y _15281_/X VGND VGND VPWR VPWR _15282_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11514_ _11513_/A _11513_/B _11513_/Y _10959_/X VGND VGND VPWR VPWR _11629_/A sky130_fd_sc_hd__o211a_1
X_14233_ _15881_/A _14250_/B VGND VGND VPWR VPWR _14233_/Y sky130_fd_sc_hd__nor2_1
X_11445_ _12346_/A _11449_/B VGND VGND VPWR VPWR _11445_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14164_ _15974_/A _14165_/B VGND VGND VPWR VPWR _14164_/X sky130_fd_sc_hd__and2_1
X_11376_ _12311_/A VGND VGND VPWR VPWR _14119_/A sky130_fd_sc_hd__buf_1
XFILLER_125_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14095_ _14095_/A _14095_/B VGND VGND VPWR VPWR _14095_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13115_ _15249_/A _13115_/B VGND VGND VPWR VPWR _13115_/Y sky130_fd_sc_hd__nand2_1
X_10327_ _10295_/X _10326_/X _10295_/X _10326_/X VGND VGND VPWR VPWR _10328_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13046_ _13032_/X _13045_/X _13032_/X _13045_/X VGND VGND VPWR VPWR _13123_/B sky130_fd_sc_hd__a2bb2o_1
X_10258_ _09268_/B _10243_/B _10243_/X _10692_/A VGND VGND VPWR VPWR _10829_/A sky130_fd_sc_hd__a22o_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10189_ _10241_/B _10151_/B _10151_/Y _10975_/A VGND VGND VPWR VPWR _10189_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14997_ _11716_/A _11723_/B _10521_/A _11716_/Y VGND VGND VPWR VPWR _14997_/X sky130_fd_sc_hd__o2bb2a_1
X_13948_ _13916_/Y _13946_/X _13947_/Y VGND VGND VPWR VPWR _13948_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13879_ _14836_/A _13980_/B _13878_/Y VGND VGND VPWR VPWR _13879_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15618_ _15616_/A _15617_/A _15616_/Y _15617_/Y _15595_/A VGND VGND VPWR VPWR _16038_/A
+ sky130_fd_sc_hd__a221o_2
X_15549_ _15497_/X _15547_/X _15579_/B VGND VGND VPWR VPWR _15549_/X sky130_fd_sc_hd__o21a_1
X_09070_ _09070_/A _09070_/B VGND VGND VPWR VPWR _09071_/B sky130_fd_sc_hd__or2_1
XFILLER_103_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09972_ _09972_/A _09972_/B VGND VGND VPWR VPWR _09972_/Y sky130_fd_sc_hd__nor2_1
X_08923_ _09292_/B VGND VGND VPWR VPWR _10228_/B sky130_fd_sc_hd__inv_2
XFILLER_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08854_ _08937_/B VGND VGND VPWR VPWR _09041_/B sky130_fd_sc_hd__inv_2
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08785_ _10012_/A VGND VGND VPWR VPWR _09470_/A sky130_fd_sc_hd__buf_1
XFILLER_29_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09406_ _09407_/A _09407_/B VGND VGND VPWR VPWR _10895_/A sky130_fd_sc_hd__and2_1
X_09337_ _08762_/A _08760_/Y _10035_/A _09336_/X VGND VGND VPWR VPWR _09337_/Y sky130_fd_sc_hd__o22ai_2
X_09268_ _09268_/A _09268_/B VGND VGND VPWR VPWR _09268_/X sky130_fd_sc_hd__or2_1
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09199_ _09199_/A VGND VGND VPWR VPWR _09199_/Y sky130_fd_sc_hd__inv_6
XFILLER_106_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11230_ _11081_/X _11229_/X _11081_/X _11229_/X VGND VGND VPWR VPWR _11231_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11161_ _11131_/X _11160_/X _11131_/X _11160_/X VGND VGND VPWR VPWR _11304_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10112_ _10112_/A _10112_/B VGND VGND VPWR VPWR _10113_/A sky130_fd_sc_hd__or2_1
X_11092_ _13901_/A _11092_/B VGND VGND VPWR VPWR _11092_/X sky130_fd_sc_hd__or2_1
XFILLER_88_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14920_ _15544_/A _14920_/B VGND VGND VPWR VPWR _14920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10043_ _10043_/A _10083_/B VGND VGND VPWR VPWR _10043_/X sky130_fd_sc_hd__and2_1
X_14851_ _14953_/A _14953_/B VGND VGND VPWR VPWR _14851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13802_ _14663_/A _13857_/B VGND VGND VPWR VPWR _13802_/Y sky130_fd_sc_hd__nor2_1
X_14782_ _14782_/A _14782_/B VGND VGND VPWR VPWR _14782_/X sky130_fd_sc_hd__and2_1
X_11994_ _11994_/A _11994_/B VGND VGND VPWR VPWR _11994_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13733_ _13695_/X _13732_/X _13695_/X _13732_/X VGND VGND VPWR VPWR _13766_/B sky130_fd_sc_hd__a2bb2o_1
X_10945_ _12162_/A VGND VGND VPWR VPWR _13702_/A sky130_fd_sc_hd__buf_1
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16452_ _16432_/X _16444_/Y _16450_/X _16451_/X VGND VGND VPWR VPWR _16472_/D sky130_fd_sc_hd__o211ai_4
X_10876_ _13078_/A _10733_/B _10733_/Y VGND VGND VPWR VPWR _10876_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13664_ _15131_/A _13629_/B _13629_/Y VGND VGND VPWR VPWR _13664_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16383_ _08230_/A _16458_/Q _08233_/A _16396_/C _16343_/A VGND VGND VPWR VPWR _16458_/D
+ sky130_fd_sc_hd__o221a_2
X_12615_ _12611_/Y _12614_/Y _12611_/A _12614_/A _12501_/A VGND VGND VPWR VPWR _14234_/B
+ sky130_fd_sc_hd__o221a_1
X_15403_ _15462_/A _15401_/X _15402_/X VGND VGND VPWR VPWR _15403_/X sky130_fd_sc_hd__o21a_1
X_15334_ _15387_/A _15332_/X _15333_/X VGND VGND VPWR VPWR _15334_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13595_ _13628_/A _13629_/B VGND VGND VPWR VPWR _13595_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12546_ _12546_/A VGND VGND VPWR VPWR _12546_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12477_ _12467_/X _12476_/Y _12467_/X _12476_/Y VGND VGND VPWR VPWR _12480_/B sky130_fd_sc_hd__a2bb2o_1
X_15265_ _15211_/A _15211_/B _15211_/Y VGND VGND VPWR VPWR _15265_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11428_ _15519_/A _11431_/B VGND VGND VPWR VPWR _12587_/A sky130_fd_sc_hd__and2_1
X_14216_ _14095_/A _14095_/B _14095_/Y VGND VGND VPWR VPWR _14216_/X sky130_fd_sc_hd__o21a_1
XANTENNA_4 _12649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15196_ _15196_/A _15196_/B VGND VGND VPWR VPWR _15196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14147_ _14066_/X _14146_/Y _14066_/X _14146_/Y VGND VGND VPWR VPWR _14148_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11359_ _08885_/X _11359_/B VGND VGND VPWR VPWR _11359_/X sky130_fd_sc_hd__and2b_1
XFILLER_112_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14078_ _14113_/A _14114_/A VGND VGND VPWR VPWR _14078_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _14591_/A _13029_/B VGND VGND VPWR VPWR _13029_/X sky130_fd_sc_hd__or2_1
XFILLER_67_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08570_ _08713_/B VGND VGND VPWR VPWR _08572_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer27 _08395_/A VGND VGND VPWR VPWR _08721_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer16 rebuffer17/X VGND VGND VPWR VPWR rebuffer16/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer49 _08375_/X VGND VGND VPWR VPWR _08455_/A1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer38 _09748_/A VGND VGND VPWR VPWR _11591_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09122_ _09122_/A VGND VGND VPWR VPWR _09122_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09053_ _08711_/Y _09052_/Y _08737_/X VGND VGND VPWR VPWR _09054_/A sky130_fd_sc_hd__o21ai_1
XFILLER_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09955_ _09955_/A _09955_/B VGND VGND VPWR VPWR _09955_/X sky130_fd_sc_hd__and2_1
XFILLER_106_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09886_/A _09886_/B VGND VGND VPWR VPWR _09887_/B sky130_fd_sc_hd__or2_1
X_08906_ _08905_/Y _08861_/X _08905_/Y _08861_/X VGND VGND VPWR VPWR _08972_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _09459_/A VGND VGND VPWR VPWR _09502_/A sky130_fd_sc_hd__buf_1
XFILLER_73_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08768_ _10132_/A VGND VGND VPWR VPWR _08768_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08699_ _08699_/A VGND VGND VPWR VPWR _08699_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_26_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10730_ _11904_/A VGND VGND VPWR VPWR _13692_/A sky130_fd_sc_hd__buf_1
X_10661_ _11023_/A _10661_/B VGND VGND VPWR VPWR _10661_/X sky130_fd_sc_hd__and2_1
XFILLER_40_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12400_ _12400_/A _12400_/B VGND VGND VPWR VPWR _12401_/B sky130_fd_sc_hd__or2_1
X_13380_ _14137_/A _13445_/B VGND VGND VPWR VPWR _13380_/Y sky130_fd_sc_hd__nor2_1
X_10592_ _10592_/A VGND VGND VPWR VPWR _10592_/Y sky130_fd_sc_hd__inv_2
X_12331_ _12331_/A _12331_/B VGND VGND VPWR VPWR _12331_/X sky130_fd_sc_hd__or2_1
X_12262_ _13712_/A _12261_/B _12261_/X _12168_/X VGND VGND VPWR VPWR _12262_/X sky130_fd_sc_hd__o22a_1
X_15050_ _15051_/A _15051_/B VGND VGND VPWR VPWR _15050_/X sky130_fd_sc_hd__and2_1
XFILLER_107_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11213_ _14023_/A _11213_/B VGND VGND VPWR VPWR _11213_/Y sky130_fd_sc_hd__nand2_1
X_14001_ _13962_/X _14000_/Y _13962_/X _14000_/Y VGND VGND VPWR VPWR _14067_/B sky130_fd_sc_hd__a2bb2o_1
X_12193_ _13719_/A _12256_/B _12192_/Y VGND VGND VPWR VPWR _12193_/Y sky130_fd_sc_hd__o21ai_1
X_11144_ _11607_/A _11144_/B VGND VGND VPWR VPWR _11145_/A sky130_fd_sc_hd__or2_1
XFILLER_1_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15952_ _15952_/A _15952_/B VGND VGND VPWR VPWR _16017_/B sky130_fd_sc_hd__or2_1
X_11075_ _12137_/A _11075_/B VGND VGND VPWR VPWR _11248_/A sky130_fd_sc_hd__and2_1
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14903_ _14046_/X _14902_/X _14046_/X _14902_/X VGND VGND VPWR VPWR _14904_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10026_ _09323_/A _08793_/B _10047_/B _10025_/X VGND VGND VPWR VPWR _10026_/X sky130_fd_sc_hd__o22a_1
X_15883_ _15886_/A _15886_/B VGND VGND VPWR VPWR _15883_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14834_ _14746_/X _14833_/Y _14764_/Y VGND VGND VPWR VPWR _14834_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14765_ _14833_/A _14833_/B _14764_/Y VGND VGND VPWR VPWR _14765_/Y sky130_fd_sc_hd__o21ai_1
X_11977_ _11945_/Y _11975_/X _11976_/Y VGND VGND VPWR VPWR _11977_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13716_ _15116_/A _13778_/B _13715_/Y VGND VGND VPWR VPWR _13716_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10928_ _10928_/A VGND VGND VPWR VPWR _10928_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16435_ _16462_/Q _16461_/Q _16464_/Q _16463_/Q VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__or4_1
X_14696_ _15343_/A _14657_/B _14657_/Y VGND VGND VPWR VPWR _14696_/Y sky130_fd_sc_hd__o21ai_1
X_10859_ _12061_/A VGND VGND VPWR VPWR _10918_/A sky130_fd_sc_hd__inv_2
X_13647_ _13538_/X _13646_/Y _13538_/X _13646_/Y VGND VGND VPWR VPWR _13648_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16366_ _16326_/A _16326_/B _16326_/Y VGND VGND VPWR VPWR _16366_/Y sky130_fd_sc_hd__o21ai_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _12847_/A _13555_/B _13556_/Y _13577_/X VGND VGND VPWR VPWR _13578_/X sky130_fd_sc_hd__o22a_1
X_16297_ _16260_/A _16326_/A _16260_/Y VGND VGND VPWR VPWR _16297_/Y sky130_fd_sc_hd__o21ai_1
X_12529_ _12634_/A _12634_/B VGND VGND VPWR VPWR _14183_/A sky130_fd_sc_hd__and2_1
X_15317_ _15337_/A _15337_/B VGND VGND VPWR VPWR _15381_/A sky130_fd_sc_hd__and2_1
XFILLER_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15248_ _15223_/X _15247_/Y _15223_/X _15247_/Y VGND VGND VPWR VPWR _15249_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15179_ _15113_/A _15113_/B _15113_/Y VGND VGND VPWR VPWR _15179_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09740_ _09740_/A _09740_/B VGND VGND VPWR VPWR _09743_/B sky130_fd_sc_hd__or2_1
.ends

