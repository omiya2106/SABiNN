VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 370.910 BY 381.630 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 365.240 104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 365.240 257.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 370.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 370.160 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 365.240 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 365.240 181.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 365.240 334.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 370.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 370.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 370.160 ;
    END
  END VPWR
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 377.630 4.050 381.630 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 201.320 370.910 201.920 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 172.760 370.910 173.360 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 340.040 370.910 340.640 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 367.240 370.910 367.840 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 257.080 370.910 257.680 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 377.630 211.050 381.630 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 377.630 61.090 381.630 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 89.800 370.910 90.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 228.520 370.910 229.120 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 377.630 286.490 381.630 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 34.040 370.910 34.640 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 377.630 248.770 381.630 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 377.630 173.330 381.630 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 377.630 229.450 381.630 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 377.630 41.770 381.630 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 6.840 370.910 7.440 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 62.600 370.910 63.200 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 377.630 304.890 381.630 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 377.630 79.490 381.630 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 377.630 267.170 381.630 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 377.630 117.210 381.630 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 377.630 192.650 381.630 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 311.480 370.910 312.080 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 377.630 361.010 381.630 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 284.280 370.910 284.880 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 377.630 154.930 381.630 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 118.360 370.910 118.960 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 377.630 342.610 381.630 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 377.630 323.290 381.630 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 377.630 97.890 381.630 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 377.630 135.610 381.630 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 377.630 23.370 381.630 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.910 145.560 370.910 146.160 ;
    END
  END wbs_dat_i[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 368.315 370.005 ;
      LAYER met1 ;
        RECT 0.070 8.540 368.375 371.580 ;
      LAYER met2 ;
        RECT 0.100 377.350 3.490 377.810 ;
        RECT 4.330 377.350 22.810 377.810 ;
        RECT 23.650 377.350 41.210 377.810 ;
        RECT 42.050 377.350 60.530 377.810 ;
        RECT 61.370 377.350 78.930 377.810 ;
        RECT 79.770 377.350 97.330 377.810 ;
        RECT 98.170 377.350 116.650 377.810 ;
        RECT 117.490 377.350 135.050 377.810 ;
        RECT 135.890 377.350 154.370 377.810 ;
        RECT 155.210 377.350 172.770 377.810 ;
        RECT 173.610 377.350 192.090 377.810 ;
        RECT 192.930 377.350 210.490 377.810 ;
        RECT 211.330 377.350 228.890 377.810 ;
        RECT 229.730 377.350 248.210 377.810 ;
        RECT 249.050 377.350 266.610 377.810 ;
        RECT 267.450 377.350 285.930 377.810 ;
        RECT 286.770 377.350 304.330 377.810 ;
        RECT 305.170 377.350 322.730 377.810 ;
        RECT 323.570 377.350 342.050 377.810 ;
        RECT 342.890 377.350 360.450 377.810 ;
        RECT 361.290 377.350 361.470 377.810 ;
        RECT 0.100 4.280 361.470 377.350 ;
        RECT 0.650 4.000 18.210 4.280 ;
        RECT 19.050 4.000 36.610 4.280 ;
        RECT 37.450 4.000 55.930 4.280 ;
        RECT 56.770 4.000 74.330 4.280 ;
        RECT 75.170 4.000 93.650 4.280 ;
        RECT 94.490 4.000 112.050 4.280 ;
        RECT 112.890 4.000 130.450 4.280 ;
        RECT 131.290 4.000 149.770 4.280 ;
        RECT 150.610 4.000 168.170 4.280 ;
        RECT 169.010 4.000 187.490 4.280 ;
        RECT 188.330 4.000 205.890 4.280 ;
        RECT 206.730 4.000 225.210 4.280 ;
        RECT 226.050 4.000 243.610 4.280 ;
        RECT 244.450 4.000 262.010 4.280 ;
        RECT 262.850 4.000 281.330 4.280 ;
        RECT 282.170 4.000 299.730 4.280 ;
        RECT 300.570 4.000 319.050 4.280 ;
        RECT 319.890 4.000 337.450 4.280 ;
        RECT 338.290 4.000 355.850 4.280 ;
        RECT 356.690 4.000 361.470 4.280 ;
      LAYER met3 ;
        RECT 3.745 368.240 366.910 370.085 ;
        RECT 3.745 366.840 366.510 368.240 ;
        RECT 3.745 361.440 366.910 366.840 ;
        RECT 4.400 360.040 366.910 361.440 ;
        RECT 3.745 341.040 366.910 360.040 ;
        RECT 3.745 339.640 366.510 341.040 ;
        RECT 3.745 334.240 366.910 339.640 ;
        RECT 4.400 332.840 366.910 334.240 ;
        RECT 3.745 312.480 366.910 332.840 ;
        RECT 3.745 311.080 366.510 312.480 ;
        RECT 3.745 305.680 366.910 311.080 ;
        RECT 4.400 304.280 366.910 305.680 ;
        RECT 3.745 285.280 366.910 304.280 ;
        RECT 3.745 283.880 366.510 285.280 ;
        RECT 3.745 278.480 366.910 283.880 ;
        RECT 4.400 277.080 366.910 278.480 ;
        RECT 3.745 258.080 366.910 277.080 ;
        RECT 3.745 256.680 366.510 258.080 ;
        RECT 3.745 249.920 366.910 256.680 ;
        RECT 4.400 248.520 366.910 249.920 ;
        RECT 3.745 229.520 366.910 248.520 ;
        RECT 3.745 228.120 366.510 229.520 ;
        RECT 3.745 222.720 366.910 228.120 ;
        RECT 4.400 221.320 366.910 222.720 ;
        RECT 3.745 202.320 366.910 221.320 ;
        RECT 3.745 200.920 366.510 202.320 ;
        RECT 3.745 194.160 366.910 200.920 ;
        RECT 4.400 192.760 366.910 194.160 ;
        RECT 3.745 173.760 366.910 192.760 ;
        RECT 3.745 172.360 366.510 173.760 ;
        RECT 3.745 166.960 366.910 172.360 ;
        RECT 4.400 165.560 366.910 166.960 ;
        RECT 3.745 146.560 366.910 165.560 ;
        RECT 3.745 145.160 366.510 146.560 ;
        RECT 3.745 139.760 366.910 145.160 ;
        RECT 4.400 138.360 366.910 139.760 ;
        RECT 3.745 119.360 366.910 138.360 ;
        RECT 3.745 117.960 366.510 119.360 ;
        RECT 3.745 111.200 366.910 117.960 ;
        RECT 4.400 109.800 366.910 111.200 ;
        RECT 3.745 90.800 366.910 109.800 ;
        RECT 3.745 89.400 366.510 90.800 ;
        RECT 3.745 84.000 366.910 89.400 ;
        RECT 4.400 82.600 366.910 84.000 ;
        RECT 3.745 63.600 366.910 82.600 ;
        RECT 3.745 62.200 366.510 63.600 ;
        RECT 3.745 55.440 366.910 62.200 ;
        RECT 4.400 54.040 366.910 55.440 ;
        RECT 3.745 35.040 366.910 54.040 ;
        RECT 3.745 33.640 366.510 35.040 ;
        RECT 3.745 28.240 366.910 33.640 ;
        RECT 4.400 26.840 366.910 28.240 ;
        RECT 3.745 7.840 366.910 26.840 ;
        RECT 3.745 6.975 366.510 7.840 ;
      LAYER met4 ;
        RECT 23.295 54.575 97.440 296.985 ;
        RECT 99.840 54.575 174.240 296.985 ;
        RECT 176.640 54.575 251.040 296.985 ;
        RECT 253.440 54.575 327.840 296.985 ;
        RECT 330.240 54.575 332.745 296.985 ;
  END
END user_project_wrapper
END LIBRARY

