magic
tech sky130A
magscale 1 2
timestamp 1637638053
<< nwell >>
rect 1066 176517 178886 177083
rect 1066 175429 178886 175995
rect 1066 174341 178886 174907
rect 1066 173253 178886 173819
rect 1066 172165 178886 172731
rect 1066 171077 178886 171643
rect 1066 169989 178886 170555
rect 1066 168901 178886 169467
rect 1066 167813 178886 168379
rect 1066 166725 178886 167291
rect 1066 165637 178886 166203
rect 1066 164549 178886 165115
rect 1066 163461 178886 164027
rect 1066 162373 178886 162939
rect 1066 161285 178886 161851
rect 1066 160197 178886 160763
rect 1066 159109 178886 159675
rect 1066 158021 178886 158587
rect 1066 156933 178886 157499
rect 1066 155845 178886 156411
rect 1066 154757 178886 155323
rect 1066 153669 178886 154235
rect 1066 152581 178886 153147
rect 1066 151493 178886 152059
rect 1066 150405 178886 150971
rect 1066 149317 178886 149883
rect 1066 148229 178886 148795
rect 1066 147141 178886 147707
rect 1066 146053 178886 146619
rect 1066 144965 178886 145531
rect 1066 143877 178886 144443
rect 1066 142789 178886 143355
rect 1066 141701 178886 142267
rect 1066 140613 178886 141179
rect 1066 139525 178886 140091
rect 1066 138437 178886 139003
rect 1066 137349 178886 137915
rect 1066 136261 178886 136827
rect 1066 135173 178886 135739
rect 1066 134085 178886 134651
rect 1066 132997 178886 133563
rect 1066 131909 178886 132475
rect 1066 130821 178886 131387
rect 1066 129733 178886 130299
rect 1066 128645 178886 129211
rect 1066 127557 178886 128123
rect 1066 126469 178886 127035
rect 1066 125381 178886 125947
rect 1066 124293 178886 124859
rect 1066 123205 178886 123771
rect 1066 122117 178886 122683
rect 1066 121029 178886 121595
rect 1066 119941 178886 120507
rect 1066 118853 178886 119419
rect 1066 117765 178886 118331
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 1104 1776 178848 177392
<< metal2 >>
rect 89994 179200 90050 180000
rect 1306 0 1362 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 9126 0 9182 800
rect 11702 0 11758 800
rect 14278 0 14334 800
rect 16946 0 17002 800
rect 19522 0 19578 800
rect 22098 0 22154 800
rect 24766 0 24822 800
rect 27342 0 27398 800
rect 29918 0 29974 800
rect 32586 0 32642 800
rect 35162 0 35218 800
rect 37830 0 37886 800
rect 40406 0 40462 800
rect 42982 0 43038 800
rect 45650 0 45706 800
rect 48226 0 48282 800
rect 50802 0 50858 800
rect 53470 0 53526 800
rect 56046 0 56102 800
rect 58622 0 58678 800
rect 61290 0 61346 800
rect 63866 0 63922 800
rect 66534 0 66590 800
rect 69110 0 69166 800
rect 71686 0 71742 800
rect 74354 0 74410 800
rect 76930 0 76986 800
rect 79506 0 79562 800
rect 82174 0 82230 800
rect 84750 0 84806 800
rect 87326 0 87382 800
rect 89994 0 90050 800
rect 92570 0 92626 800
rect 95238 0 95294 800
rect 97814 0 97870 800
rect 100390 0 100446 800
rect 103058 0 103114 800
rect 105634 0 105690 800
rect 108210 0 108266 800
rect 110878 0 110934 800
rect 113454 0 113510 800
rect 116030 0 116086 800
rect 118698 0 118754 800
rect 121274 0 121330 800
rect 123942 0 123998 800
rect 126518 0 126574 800
rect 129094 0 129150 800
rect 131762 0 131818 800
rect 134338 0 134394 800
rect 136914 0 136970 800
rect 139582 0 139638 800
rect 142158 0 142214 800
rect 144734 0 144790 800
rect 147402 0 147458 800
rect 149978 0 150034 800
rect 152646 0 152702 800
rect 155222 0 155278 800
rect 157798 0 157854 800
rect 160466 0 160522 800
rect 163042 0 163098 800
rect 165618 0 165674 800
rect 168286 0 168342 800
rect 170862 0 170918 800
rect 173438 0 173494 800
rect 176106 0 176162 800
rect 178682 0 178738 800
<< obsm2 >>
rect 1306 856 178736 177392
rect 1418 734 3826 856
rect 3994 734 6402 856
rect 6570 734 9070 856
rect 9238 734 11646 856
rect 11814 734 14222 856
rect 14390 734 16890 856
rect 17058 734 19466 856
rect 19634 734 22042 856
rect 22210 734 24710 856
rect 24878 734 27286 856
rect 27454 734 29862 856
rect 30030 734 32530 856
rect 32698 734 35106 856
rect 35274 734 37774 856
rect 37942 734 40350 856
rect 40518 734 42926 856
rect 43094 734 45594 856
rect 45762 734 48170 856
rect 48338 734 50746 856
rect 50914 734 53414 856
rect 53582 734 55990 856
rect 56158 734 58566 856
rect 58734 734 61234 856
rect 61402 734 63810 856
rect 63978 734 66478 856
rect 66646 734 69054 856
rect 69222 734 71630 856
rect 71798 734 74298 856
rect 74466 734 76874 856
rect 77042 734 79450 856
rect 79618 734 82118 856
rect 82286 734 84694 856
rect 84862 734 87270 856
rect 87438 734 89938 856
rect 90106 734 92514 856
rect 92682 734 95182 856
rect 95350 734 97758 856
rect 97926 734 100334 856
rect 100502 734 103002 856
rect 103170 734 105578 856
rect 105746 734 108154 856
rect 108322 734 110822 856
rect 110990 734 113398 856
rect 113566 734 115974 856
rect 116142 734 118642 856
rect 118810 734 121218 856
rect 121386 734 123886 856
rect 124054 734 126462 856
rect 126630 734 129038 856
rect 129206 734 131706 856
rect 131874 734 134282 856
rect 134450 734 136858 856
rect 137026 734 139526 856
rect 139694 734 142102 856
rect 142270 734 144678 856
rect 144846 734 147346 856
rect 147514 734 149922 856
rect 150090 734 152590 856
rect 152758 734 155166 856
rect 155334 734 157742 856
rect 157910 734 160410 856
rect 160578 734 162986 856
rect 163154 734 165562 856
rect 165730 734 168230 856
rect 168398 734 170806 856
rect 170974 734 173382 856
rect 173550 734 176050 856
rect 176218 734 178626 856
<< metal3 >>
rect 179200 90040 180000 90160
<< obsm3 >>
rect 1301 90240 179200 177377
rect 1301 89960 179120 90240
rect 1301 2143 179200 89960
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< obsm4 >>
rect 8155 10099 19488 59533
rect 19968 10099 34848 59533
rect 35328 10099 48149 59533
<< labels >>
rlabel metal2 s 89994 179200 90050 180000 6 user_clock2
port 1 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 user_irq[0]
port 2 nsew signal output
rlabel metal3 s 179200 90040 180000 90160 6 user_irq[1]
port 3 nsew signal output
rlabel metal2 s 178682 0 178738 800 6 user_irq[2]
port 4 nsew signal output
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 5 nsew power input
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 5 nsew power input
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 5 nsew power input
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 5 nsew power input
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 5 nsew power input
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 5 nsew power input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 6 nsew ground input
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 6 nsew ground input
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 6 nsew ground input
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 6 nsew ground input
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 6 nsew ground input
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 6 nsew ground input
rlabel metal2 s 1306 0 1362 800 6 wb_clk_i
port 7 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wb_rst_i
port 8 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_ack_o
port 9 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[0]
port 10 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 wbs_adr_i[10]
port 11 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 wbs_adr_i[11]
port 12 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 wbs_adr_i[12]
port 13 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_adr_i[13]
port 14 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_adr_i[14]
port 15 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 wbs_adr_i[15]
port 16 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 wbs_adr_i[16]
port 17 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 wbs_adr_i[17]
port 18 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 wbs_adr_i[18]
port 19 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 wbs_adr_i[19]
port 20 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[1]
port 21 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 wbs_adr_i[20]
port 22 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 wbs_adr_i[21]
port 23 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 wbs_adr_i[22]
port 24 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 wbs_adr_i[23]
port 25 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 wbs_adr_i[24]
port 26 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 wbs_adr_i[25]
port 27 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 wbs_adr_i[26]
port 28 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 wbs_adr_i[27]
port 29 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 wbs_adr_i[28]
port 30 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 wbs_adr_i[29]
port 31 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[2]
port 32 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 wbs_adr_i[30]
port 33 nsew signal input
rlabel metal2 s 170862 0 170918 800 6 wbs_adr_i[31]
port 34 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[3]
port 35 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[4]
port 36 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[5]
port 37 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_adr_i[6]
port 38 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 wbs_adr_i[7]
port 39 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_adr_i[8]
port 40 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_adr_i[9]
port 41 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[0]
port 42 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 wbs_dat_i[10]
port 43 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 wbs_dat_i[11]
port 44 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 wbs_dat_i[12]
port 45 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 wbs_dat_i[13]
port 46 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_i[14]
port 47 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_i[15]
port 48 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 wbs_dat_i[16]
port 49 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_dat_i[17]
port 50 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 wbs_dat_i[18]
port 51 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 wbs_dat_i[19]
port 52 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[1]
port 53 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 wbs_dat_i[20]
port 54 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 wbs_dat_i[21]
port 55 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_i[22]
port 56 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 wbs_dat_i[23]
port 57 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 wbs_dat_i[24]
port 58 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 wbs_dat_i[25]
port 59 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 wbs_dat_i[26]
port 60 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 wbs_dat_i[27]
port 61 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 wbs_dat_i[28]
port 62 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 wbs_dat_i[29]
port 63 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[2]
port 64 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 wbs_dat_i[30]
port 65 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 wbs_dat_i[31]
port 66 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_i[3]
port 67 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_i[4]
port 68 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[5]
port 69 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_i[6]
port 70 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_i[7]
port 71 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_i[8]
port 72 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_i[9]
port 73 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 180000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 27340942
string GDS_START 675022
<< end >>

